//: version "1.8.7"

module main;    //: root_module
wire w6;    //: /sn:0 {0}(291,237)(476,237)(476,251){1}
wire w16;    //: /sn:0 {0}(292,527)(473,527)(473,543){1}
wire w14;    //: /sn:0 {0}(409,450)(394,450)(394,520)(520,520)(520,603)(510,603){1}
wire w19;    //: /sn:0 /dp:1 {0}(458,660)(458,667)(580,667)(580,612)(647,612)(647,551)(704,551){1}
wire w15;    //: /sn:0 {0}(197,533)(425,533)(425,543){1}
wire w4;    //: /sn:0 {0}(409,163)(396,163)(396,230)(521,230)(521,305)(511,305){1}
wire w3;    //: /sn:0 {0}(460,208)(460,216)(591,216)(591,581)(704,581){1}
wire w0;    //: /sn:0 {0}(197,97)(427,97)(427,108){1}
wire [3:0] w21;    //: /sn:0 {0}(287,56)(287,84){1}
//: {2}(287,85)(287,236){3}
//: {4}(287,237)(287,377){5}
//: {6}(287,378)(287,452)(288,452)(288,526){7}
//: {8}(288,527)(288,620){9}
wire [3:0] w20;    //: /sn:0 {0}(190,57)(190,75)(193,75)(193,96){1}
//: {2}(193,97)(193,243){3}
//: {4}(193,244)(193,388){5}
//: {6}(193,389)(193,532){7}
//: {8}(193,533)(193,621){9}
wire w1;    //: /sn:0 {0}(291,85)(474,85)(474,108){1}
wire w8;    //: /sn:0 {0}(456,351)(456,361)(605,361)(605,571)(704,571){1}
wire [3:0] w17;    //: /sn:0 {0}(710,566)(852,566)(852,520){1}
wire w22;    //: /sn:0 {0}(580,96)(590,96)(590,165)(514,165){1}
wire w2;    //: /sn:0 {0}(355,575)(355,604)(406,604){1}
wire w11;    //: /sn:0 {0}(291,378)(484,378)(484,396){1}
wire w10;    //: /sn:0 {0}(197,389)(443,389)(443,396){1}
wire w13;    //: /sn:0 /dp:1 {0}(459,502)(459,510)(560,510)(560,561)(704,561){1}
wire w5;    //: /sn:0 {0}(197,244)(432,244)(432,251){1}
wire w9;    //: /sn:0 {0}(404,302)(394,302)(394,372)(523,372)(523,446)(513,446){1}
//: enddecls

  tran g8(.Z(w15), .I(w20[3]));   //: @(191,533) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: dip g4 (w20) @(190,47) /sn:0 /w:[ 0 ] /st:0
  tran g13(.Z(w16), .I(w21[3]));   //: @(286,527) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  FA g3 (.b(w16), .a(w15), .Cin(w14), .Cout(w2), .s(w19));   //: @(407, 544) /sz:(102, 115) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  FA g2 (.b(w11), .a(w10), .Cin(w9), .Cout(w14), .s(w13));   //: @(410, 397) /sz:(102, 104) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FA g1 (.b(w6), .a(w5), .Cin(w4), .Cout(w9), .s(w8));   //: @(405, 252) /sz:(105, 98) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  concat g16 (.I0(w3), .I1(w8), .I2(w13), .I3(w19), .Z(w17));   //: @(709,566) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  tran g11(.Z(w6), .I(w21[1]));   //: @(285,237) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  tran g10(.Z(w1), .I(w21[0]));   //: @(285,85) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  tran g6(.Z(w5), .I(w20[1]));   //: @(191,244) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: dip g9 (w21) @(287,46) /sn:0 /w:[ 0 ] /st:0
  tran g7(.Z(w10), .I(w20[2]));   //: @(191,389) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  led g15 (.I(w2));   //: @(355,568) /sn:0 /w:[ 0 ] /type:0
  led g17 (.I(w17));   //: @(852,513) /sn:0 /w:[ 1 ] /type:3
  //: switch g14 (w22) @(563,96) /sn:0 /w:[ 0 ] /st:0
  tran g5(.Z(w0), .I(w20[0]));   //: @(191,97) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  FA g0 (.b(w1), .a(w0), .Cin(w22), .Cout(w4), .s(w3));   //: @(410, 109) /sz:(103, 98) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  tran g12(.Z(w11), .I(w21[2]));   //: @(285,378) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1

endmodule

module FA(s, b, Cout, Cin, a);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(428,286)(453,286){1}
//: {2}(457,286)(486,286)(486,278)(494,278){3}
//: {4}(455,288)(455,353)(581,353){5}
output Cout;    //: /sn:0 {0}(695,338)(676,338){1}
input Cin;    //: /sn:0 {0}(427,306)(573,306){1}
//: {2}(575,304)(575,281)(585,281){3}
//: {4}(575,308)(575,318)(582,318){5}
output s;    //: /sn:0 /dp:1 {0}(606,279)(695,279){1}
input a;    //: /sn:0 {0}(426,273)(444,273){1}
//: {2}(448,273)(494,273){3}
//: {4}(446,275)(446,358)(581,358){5}
wire w8;    //: /sn:0 {0}(603,321)(645,321)(645,335)(655,335){1}
wire w11;    //: /sn:0 {0}(602,356)(645,356)(645,340)(655,340){1}
wire w2;    //: /sn:0 {0}(515,276)(525,276){1}
//: {2}(529,276)(585,276){3}
//: {4}(527,278)(527,323)(582,323){5}
//: enddecls

  //: output g8 (s) @(692,279) /sn:0 /w:[ 1 ]
  or g4 (.I0(w8), .I1(w11), .Z(Cout));   //: @(666,338) /sn:0 /delay:" 3" /w:[ 1 1 1 ]
  //: joint g13 (Cin) @(575, 306) /w:[ -1 2 1 4 ]
  and g3 (.I0(b), .I1(a), .Z(w11));   //: @(592,356) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  and g2 (.I0(Cin), .I1(w2), .Z(w8));   //: @(593,321) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  xor g1 (.I0(w2), .I1(Cin), .Z(s));   //: @(596,279) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: joint g11 (b) @(455, 286) /w:[ 2 -1 1 4 ]
  //: joint g10 (a) @(446, 273) /w:[ 2 -1 1 4 ]
  //: input g6 (b) @(426,286) /sn:0 /w:[ 0 ]
  //: output g9 (Cout) @(692,338) /sn:0 /w:[ 0 ]
  //: input g7 (Cin) @(425,306) /sn:0 /w:[ 0 ]
  //: input g5 (a) @(424,273) /sn:0 /w:[ 0 ]
  xor g0 (.I0(a), .I1(b), .Z(w2));   //: @(505,276) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: joint g12 (w2) @(527, 276) /w:[ 2 -1 1 4 ]

endmodule
