//: version "1.8.7"

module main;    //: root_module
wire w6;    //: /sn:0 {0}(272,355)(272,365)(290,365)(290,326){1}
wire w7;    //: /sn:0 {0}(333,354)(333,364)(356,364)(356,326){1}
wire w4;    //: /sn:0 {0}(351,91)(360,91)(360,131){1}
wire w3;    //: /sn:0 {0}(279,92)(288,92)(288,131){1}
wire w8;    //: /sn:0 {0}(402,353)(402,363)(425,363)(425,326){1}
wire w5;    //: /sn:0 {0}(415,92)(425,92)(425,131){1}
//: enddecls

  //: switch g4 (w3) @(262,92) /sn:0 /w:[ 0 ] /st:0
  led g3 (.I(w8));   //: @(402,346) /sn:0 /w:[ 0 ] /type:0
  led g2 (.I(w7));   //: @(333,347) /sn:0 /w:[ 0 ] /type:0
  led g1 (.I(w6));   //: @(272,348) /sn:0 /w:[ 0 ] /type:0
  //: switch g6 (w5) @(398,92) /sn:0 /w:[ 0 ] /st:0
  //: switch g5 (w4) @(334,91) /sn:0 /w:[ 0 ] /st:0
  PFA g0 (.c(w5), .b(w4), .a(w3), .g(w6), .p(w7), .s(w8));   //: @(256, 132) /sz:(216, 193) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<1 Bo1<1 Bo2<1 ]

endmodule

module PFA(s, b, g, a, c, p);
//: interface  /sz:(40, 40) /bd:[ ]
output p;    //: /sn:0 /dp:1 {0}(491,244)(543,244){1}
input b;    //: /sn:0 {0}(478,288)(337,288)(337,248){1}
//: {2}(339,246)(470,246){3}
//: {4}(337,244)(337,186){5}
//: {6}(339,184)(375,184)(375,174)(383,174){7}
//: {8}(335,184)(322,184){9}
output s;    //: /sn:0 /dp:1 {0}(497,205)(543,205){1}
input a;    //: /sn:0 /dp:9 {0}(478,283)(351,283)(351,243){1}
//: {2}(353,241)(470,241){3}
//: {4}(351,239)(351,171){5}
//: {6}(353,169)(383,169){7}
//: {8}(349,169)(322,169){9}
output g;    //: /sn:0 /dp:1 {0}(499,286)(521,286)(521,284)(543,284){1}
input c;    //: /sn:0 {0}(322,207)(476,207){1}
wire w2;    //: /sn:0 {0}(404,172)(468,172)(468,202)(476,202){1}
//: enddecls

  //: output g4 (s) @(540,205) /sn:0 /w:[ 1 ]
  //: input g8 (b) @(320,184) /sn:0 /w:[ 9 ]
  and g3 (.I0(a), .I1(b), .Z(g));   //: @(489,286) /sn:0 /delay:" 3" /w:[ 0 0 0 ]
  //: joint g13 (a) @(351, 241) /w:[ 2 4 -1 1 ]
  or g2 (.I0(a), .I1(b), .Z(p));   //: @(481,244) /sn:0 /delay:" 3" /w:[ 3 3 0 ]
  xor g1 (.I0(w2), .I1(c), .Z(s));   //: @(487,205) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  //: joint g11 (b) @(337, 246) /w:[ 2 4 -1 1 ]
  //: joint g10 (a) @(351, 169) /w:[ 6 -1 8 5 ]
  //: output g6 (g) @(540,284) /sn:0 /w:[ 1 ]
  //: input g7 (a) @(320,169) /sn:0 /w:[ 9 ]
  //: input g9 (c) @(320,207) /sn:0 /w:[ 0 ]
  //: output g5 (p) @(540,244) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(w2));   //: @(394,172) /sn:0 /delay:" 4" /w:[ 7 7 0 ]
  //: joint g12 (b) @(337, 184) /w:[ 6 -1 8 5 ]

endmodule
