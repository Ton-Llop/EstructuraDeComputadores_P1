//: version "1.8.7"

module restador(Cout, b, a, S);
//: interface  /sz:(40, 40) /bd:[ ]
input [15:0] b;    //: /sn:0 {0}(199,20)(199,58){1}
supply1 w0;    //: /sn:0 {0}(272,102)(272,133)(211,133){1}
output Cout;    //: /sn:0 {0}(8,116)(131,116)(131,136)(169,136){1}
input [15:0] a;    //: /sn:0 {0}(143,83)(179,83)(179,107){1}
output [15:0] S;    //: /sn:0 {0}(190,149)(190,174)(218,174){1}
wire [15:0] w5;    //: /sn:0 {0}(199,74)(199,107){1}
//: enddecls

  //: output g4 (Cout) @(11,116) /sn:0 /R:2 /w:[ 0 ]
  not g3 (.I(b), .Z(w5));   //: @(199,64) /sn:0 /R:3 /w:[ 1 0 ]
  //: input g2 (b) @(199,18) /sn:0 /R:3 /w:[ 0 ]
  //: input g1 (a) @(141,83) /sn:0 /w:[ 0 ]
  //: output g6 (S) @(215,174) /sn:0 /w:[ 1 ]
  //: supply1 g5 (w0) @(283,102) /sn:0 /w:[ 0 ]
  CPA16B g0 (.b(w5), .a(a), .Cin(w0), .Cout(Cout), .S(S));   //: @(170, 108) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]

endmodule

module CPA(b, a, Cin, s, Cout);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] b;    //: /sn:0 {0}(72,53)(86,53)(86,143)(305,143){1}
//: {2}(306,143)(515,143){3}
//: {4}(516,143)(717,143){5}
//: {6}(718,143)(922,143){7}
//: {8}(923,143)(967,143){9}
output Cout;    //: /sn:0 {0}(971,250)(1035,250){1}
input Cin;    //: /sn:0 {0}(104,237)(217,237)(217,261)(227,261){1}
output [3:0] s;    //: /sn:0 /dp:1 {0}(983,407)(1099,407)(1099,387)(1103,387){1}
input [3:0] a;    //: /sn:0 {0}(135,60)(143,60)(143,124)(255,124){1}
//: {2}(256,124)(462,124){3}
//: {4}(463,124)(677,124){5}
//: {6}(678,124)(871,124){7}
//: {8}(872,124)(1006,124){9}
wire w6;    //: /sn:0 {0}(516,147)(516,185){1}
wire w7;    //: /sn:0 {0}(577,254)(632,254)(632,261)(642,261){1}
wire w16;    //: /sn:0 {0}(923,147)(923,183){1}
wire w15;    //: /sn:0 {0}(872,128)(872,183){1}
wire w3;    //: /sn:0 {0}(351,256)(411,256)(411,257)(421,257){1}
wire w0;    //: /sn:0 {0}(256,128)(256,187){1}
wire w1;    //: /sn:0 {0}(306,147)(306,155)(307,155)(307,187){1}
wire w18;    //: /sn:0 /dp:1 {0}(907,328)(907,392)(977,392){1}
wire w8;    //: /sn:0 {0}(498,325)(498,412)(977,412){1}
wire w12;    //: /sn:0 {0}(767,256)(843,256){1}
wire w11;    //: /sn:0 {0}(718,147)(718,185){1}
wire w2;    //: /sn:0 {0}(290,324)(290,422)(977,422){1}
wire w10;    //: /sn:0 {0}(678,128)(678,185){1}
wire w13;    //: /sn:0 /dp:1 {0}(705,329)(705,402)(977,402){1}
wire w5;    //: /sn:0 {0}(463,128)(463,154)(462,154)(462,185){1}
//: enddecls

  //: input g8 (b) @(70,53) /sn:0 /w:[ 0 ]
  //: input g4 (a) @(133,60) /sn:0 /w:[ 0 ]
  //: input g13 (Cin) @(102,237) /sn:0 /w:[ 0 ]
  FA g3 (.b(w16), .a(w15), .Cin(w12), .s(w18), .Cout(Cout));   //: @(844, 184) /sz:(126, 143) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  FA g2 (.b(w11), .a(w10), .Cin(w7), .s(w13), .Cout(w12));   //: @(643, 186) /sz:(123, 142) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  FA g1 (.b(w6), .a(w5), .Cin(w3), .s(w8), .Cout(w7));   //: @(422, 186) /sz:(154, 138) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  //: output g16 (s) @(1100,387) /sn:0 /w:[ 1 ]
  tran g11(.Z(w11), .I(b[2]));   //: @(718,141) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g10(.Z(w6), .I(b[1]));   //: @(516,141) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g6(.Z(w5), .I(a[1]));   //: @(463,122) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g9(.Z(w1), .I(b[0]));   //: @(306,141) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g7(.Z(w10), .I(a[2]));   //: @(678,122) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  concat g15 (.I0(w2), .I1(w8), .I2(w13), .I3(w18), .Z(s));   //: @(982,407) /sn:0 /w:[ 1 1 1 1 0 ] /dr:0
  //: output g14 (Cout) @(1032,250) /sn:0 /w:[ 1 ]
  tran g5(.Z(w0), .I(a[0]));   //: @(256,122) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  FA g0 (.b(w1), .a(w0), .Cin(Cin), .s(w2), .Cout(w3));   //: @(228, 188) /sz:(122, 135) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  tran g12(.Z(w16), .I(b[3]));   //: @(923,141) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran D4(.Z(w15), .I(a[3]));   //: @(872,122) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1

endmodule

module CPA16B(a, S, b, Cout, Cin);
//: interface  /sz:(40, 40) /bd:[ ]
input [15:0] b;    //: /sn:0 {0}(-11,92)(46,92)(46,119)(315,119){1}
//: {2}(316,119)(568,119){3}
//: {4}(569,119)(809,119){5}
//: {6}(810,119)(1049,119){7}
//: {8}(1050,119)(1115,119){9}
output Cout;    //: /sn:0 {0}(1270,287)(1131,287)(1131,251)(1121,251){1}
input Cin;    //: /sn:0 /dp:1 {0}(197,253)(144,253)(144,231)(108,231){1}
input [15:0] a;    //: /sn:0 {0}(-21,52)(101,52)(101,97)(239,97){1}
//: {2}(240,97)(372,97)(372,99)(504,99){3}
//: {4}(505,99)(760,99){5}
//: {6}(761,99)(981,99){7}
//: {8}(982,99)(1114,99){9}
output [15:0] S;    //: /sn:0 /dp:1 {0}(1304,487)(1291,487)(1291,498)(1197,498){1}
wire [3:0] w6;    //: /sn:0 {0}(569,123)(569,131)(570,131)(570,151){1}
wire w7;    //: /sn:0 {0}(626,255)(693,255){1}
wire [3:0] w16;    //: /sn:0 {0}(1050,123)(1050,153){1}
wire [3:0] w14;    //: /sn:0 {0}(779,342)(779,493)(1191,493){1}
wire [3:0] w15;    //: /sn:0 {0}(982,103)(982,153){1}
wire [3:0] w4;    //: /sn:0 /dp:1 {0}(1191,513)(1130,513)(1130,527)(283,527)(283,345){1}
wire w3;    //: /sn:0 {0}(374,251)(412,251)(412,253)(452,253){1}
wire [3:0] w0;    //: /sn:0 {0}(240,101)(240,124)(239,124)(239,149){1}
wire [3:0] w24;    //: /sn:0 {0}(1191,483)(1107,483)(1107,467)(1027,467)(1027,338){1}
wire [3:0] w1;    //: /sn:0 {0}(316,123)(316,135)(315,135)(315,149){1}
wire [3:0] w11;    //: /sn:0 {0}(810,123)(810,154){1}
wire [3:0] w10;    //: /sn:0 {0}(761,103)(761,154){1}
wire w13;    //: /sn:0 {0}(873,253)(940,253){1}
wire [3:0] w5;    //: /sn:0 {0}(505,103)(505,151){1}
wire [3:0] w9;    //: /sn:0 {0}(534,347)(534,503)(1191,503){1}
//: enddecls

  tran g8(.Z(w15), .I(a[15:12]));   //: @(982,97) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: input g4 (a) @(-23,52) /sn:0 /w:[ 0 ]
  CPA g3 (.b(w16), .a(w15), .Cin(w13), .s(w24), .Cout(Cout));   //: @(941, 154) /sz:(179, 183) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<1 Ro0<1 ]
  tran g13(.Z(w16), .I(b[15:12]));   //: @(1050,117) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  CPA g2 (.b(w11), .a(w10), .Cin(w7), .s(w14), .Cout(w13));   //: @(694, 155) /sz:(178, 186) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  CPA g1 (.b(w6), .a(w5), .Cin(w3), .s(w9), .Cout(w7));   //: @(453, 152) /sz:(172, 194) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  tran g11(.Z(w6), .I(b[7:4]));   //: @(569,117) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: output g16 (S) @(1301,487) /sn:0 /w:[ 0 ]
  tran g10(.Z(w1), .I(b[3:0]));   //: @(316,117) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g6(.Z(w5), .I(a[7:4]));   //: @(505,97) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g7(.Z(w10), .I(a[11:8]));   //: @(761,97) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: input g9 (b) @(-13,92) /sn:0 /w:[ 0 ]
  concat g15 (.I0(w4), .I1(w9), .I2(w14), .I3(w24), .Z(S));   //: @(1196,498) /sn:0 /w:[ 0 1 1 0 1 ] /dr:0
  //: output g17 (Cout) @(1267,287) /sn:0 /w:[ 0 ]
  tran g5(.Z(w0), .I(a[3:0]));   //: @(240,95) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g14 (Cin) @(106,231) /sn:0 /w:[ 1 ]
  CPA g0 (.b(w1), .a(w0), .Cin(Cin), .s(w4), .Cout(w3));   //: @(198, 150) /sz:(175, 194) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>0 Bo0<1 Ro0<0 ]
  tran g12(.Z(w11), .I(b[11:8]));   //: @(810,117) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w4;    //: /sn:0 /dp:1 {0}(339,135)(339,192)(382,192)(382,202){1}
wire [15:0] w0;    //: /sn:0 /dp:1 {0}(435,131)(435,193)(403,193)(403,202){1}
wire [15:0] w1;    //: /sn:0 {0}(543,271)(543,281)(382,281)(382,244){1}
wire w2;    //: /sn:0 {0}(418,226)(471,226){1}
//: enddecls

  led g4 (.I(w1));   //: @(543,264) /sn:0 /w:[ 0 ] /type:2
  led g3 (.I(w2));   //: @(478,226) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: dip g2 (w0) @(435,121) /sn:0 /w:[ 0 ] /st:0
  //: dip g1 (w4) @(339,125) /sn:0 /w:[ 0 ] /st:0
  restador g0 (.b(w0), .a(w4), .S(w1), .Cout(w2));   //: @(377, 203) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 Ro0<0 ]

endmodule

module FA(s, b, Cin, Cout, a);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(428,286)(453,286){1}
//: {2}(457,286)(486,286)(486,278)(494,278){3}
//: {4}(455,288)(455,353)(581,353){5}
output Cout;    //: /sn:0 {0}(695,338)(676,338){1}
input Cin;    //: /sn:0 {0}(427,306)(573,306){1}
//: {2}(575,304)(575,281)(585,281){3}
//: {4}(575,308)(575,318)(582,318){5}
output s;    //: /sn:0 /dp:1 {0}(606,279)(695,279){1}
input a;    //: /sn:0 {0}(426,273)(444,273){1}
//: {2}(448,273)(494,273){3}
//: {4}(446,275)(446,358)(581,358){5}
wire w8;    //: /sn:0 {0}(603,321)(645,321)(645,335)(655,335){1}
wire w2;    //: /sn:0 {0}(515,276)(525,276){1}
//: {2}(529,276)(585,276){3}
//: {4}(527,278)(527,323)(582,323){5}
wire w11;    //: /sn:0 {0}(602,356)(645,356)(645,340)(655,340){1}
//: enddecls

  or g4 (.I0(w8), .I1(w11), .Z(Cout));   //: @(666,338) /sn:0 /delay:" 3" /w:[ 1 1 1 ]
  //: output g8 (s) @(692,279) /sn:0 /w:[ 1 ]
  and g3 (.I0(b), .I1(a), .Z(w11));   //: @(592,356) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: joint g13 (Cin) @(575, 306) /w:[ -1 2 1 4 ]
  and g2 (.I0(Cin), .I1(w2), .Z(w8));   //: @(593,321) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  xor g1 (.I0(w2), .I1(Cin), .Z(s));   //: @(596,279) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: joint g11 (b) @(455, 286) /w:[ 2 -1 1 4 ]
  //: joint g10 (a) @(446, 273) /w:[ 2 -1 1 4 ]
  //: input g6 (b) @(426,286) /sn:0 /w:[ 0 ]
  //: input g7 (Cin) @(425,306) /sn:0 /w:[ 0 ]
  //: output g9 (Cout) @(692,338) /sn:0 /w:[ 0 ]
  //: input g5 (a) @(424,273) /sn:0 /w:[ 0 ]
  xor g0 (.I0(a), .I1(b), .Z(w2));   //: @(505,276) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: joint g12 (w2) @(527, 276) /w:[ 2 -1 1 4 ]

endmodule
