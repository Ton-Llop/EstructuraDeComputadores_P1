//: version "1.8.7"

module FAalternativa(Cout, b, Cin, s, a);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(233,117)(278,117){1}
//: {2}(282,117)(354,117){3}
//: {4}(280,119)(280,212){5}
//: {6}(282,214)(359,214){7}
//: {8}(280,216)(280,256)(358,256){9}
output Cout;    //: /sn:0 /dp:1 {0}(478,212)(515,212){1}
input Cin;    //: /sn:0 {0}(232,139)(255,139){1}
//: {2}(259,139)(319,139){3}
//: {4}(323,139)(346,139)(346,122)(354,122){5}
//: {6}(321,141)(321,173)(357,173){7}
//: {8}(257,141)(257,261)(358,261){9}
output s;    //: /sn:0 /dp:1 {0}(375,117)(384,117)(384,127)(393,127)(393,117){1}
//: {2}(395,115)(434,115)(434,115)(451,115){3}
//: {4}(391,115)(383,115){5}
input a;    //: /sn:0 {0}(235,106)(250,106){1}
//: {2}(254,106)(346,106)(346,112)(354,112){3}
//: {4}(252,104)(252,93)(267,93)(267,209)(359,209){5}
//: {6}(252,108)(252,178)(357,178){7}
wire w6;    //: /sn:0 {0}(378,176)(445,176)(445,207)(457,207){1}
wire w12;    //: /sn:0 {0}(379,259)(446,259)(446,217)(457,217){1}
wire w9;    //: /sn:0 {0}(380,212)(457,212){1}
//: enddecls

  //: output g8 (Cout) @(512,212) /sn:0 /w:[ 1 ]
  or g4 (.I0(w6), .I1(w9), .I2(w12), .Z(Cout));   //: @(468,212) /sn:0 /delay:" 3" /w:[ 1 1 1 0 ]
  and g3 (.I0(b), .I1(Cin), .Z(w12));   //: @(369,259) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: joint g13 (b) @(280, 117) /w:[ 2 -1 1 4 ]
  and g2 (.I0(a), .I1(b), .Z(w9));   //: @(370,212) /sn:0 /delay:" 3" /w:[ 5 7 0 ]
  and g1 (.I0(Cin), .I1(a), .Z(w6));   //: @(368,176) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: joint g11 (Cin) @(321, 139) /w:[ 4 -1 3 6 ]
  //: joint g10 (s) @(393, 115) /w:[ 2 -1 4 1 ]
  //: input g6 (b) @(231,117) /sn:0 /w:[ 0 ]
  //: input g7 (Cin) @(230,139) /sn:0 /w:[ 0 ]
  //: output g9 (s) @(448,115) /sn:0 /w:[ 3 ]
  //: joint g15 (Cin) @(257, 139) /w:[ 2 -1 1 8 ]
  //: input g5 (a) @(233,106) /sn:0 /w:[ 0 ]
  //: joint g14 (b) @(280, 214) /w:[ 6 5 -1 8 ]
  xor g0 (.I0(a), .I1(b), .I2(Cin), .Z(s));   //: @(365,117) /sn:0 /delay:" 4" /w:[ 3 3 5 0 ]
  //: joint g12 (a) @(252, 106) /w:[ 2 4 1 6 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(396,446)(396,466)(429,466)(429,406){1}
wire w0;    //: /sn:0 {0}(449,57)(472,57)(472,123){1}
wire w3;    //: /sn:0 {0}(317,59)(333,59)(333,123){1}
wire w1;    //: /sn:0 {0}(672,221)(682,221)(682,265)(602,265){1}
wire w5;    //: /sn:0 {0}(218,236)(218,266)(253,266){1}
//: enddecls

  //: switch g4 (w0) @(432,57) /sn:0 /w:[ 0 ] /st:0
  //: switch g3 (w3) @(300,59) /sn:0 /w:[ 0 ] /st:0
  led g2 (.I(w4));   //: @(396,439) /sn:0 /w:[ 0 ] /type:0
  led g1 (.I(w5));   //: @(218,229) /sn:0 /w:[ 0 ] /type:0
  //: switch g5 (w1) @(655,221) /sn:0 /w:[ 0 ] /st:0
  FAalternativa g0 (.b(w0), .a(w3), .Cin(w1), .Cout(w5), .s(w4));   //: @(254, 124) /sz:(347, 281) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]

endmodule
