//: version "1.8.7"

module FAalterniva(s, b, Cout, Cin, a);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(269,176)(330,176){1}
//: {2}(334,176)(396,176){3}
//: {4}(332,178)(332,293){5}
//: {6}(334,295)(391,295){7}
//: {8}(332,297)(332,329)(391,329){9}
output Cout;    //: /sn:0 /dp:1 {0}(525,293)(563,293){1}
input Cin;    //: /sn:0 {0}(268,201)(284,201){1}
//: {2}(288,201)(348,201){3}
//: {4}(352,201)(388,201)(388,181)(396,181){5}
//: {6}(350,203)(350,245)(390,245){7}
//: {8}(286,203)(286,334)(391,334){9}
output s;    //: /sn:0 /dp:1 {0}(417,176)(524,176){1}
input a;    //: /sn:0 {0}(268,154)(299,154){1}
//: {2}(303,154)(388,154)(388,171)(396,171){3}
//: {4}(301,152)(301,142)(316,142)(316,290)(391,290){5}
//: {6}(301,156)(301,250)(390,250){7}
wire w8;    //: /sn:0 {0}(412,293)(504,293){1}
wire w11;    //: /sn:0 {0}(412,332)(492,332)(492,298)(504,298){1}
wire w5;    //: /sn:0 {0}(411,248)(494,248)(494,288)(504,288){1}
//: enddecls

  //: output g8 (s) @(521,176) /sn:0 /w:[ 1 ]
  or g4 (.I0(w5), .I1(w8), .I2(w11), .Z(Cout));   //: @(515,293) /sn:0 /delay:" 3" /w:[ 1 1 1 0 ]
  //: joint g13 (Cin) @(350, 201) /w:[ 4 -1 3 6 ]
  and g3 (.I0(b), .I1(Cin), .Z(w11));   //: @(402,332) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  and g2 (.I0(a), .I1(b), .Z(w8));   //: @(402,293) /sn:0 /delay:" 3" /w:[ 5 7 0 ]
  and g1 (.I0(Cin), .I1(a), .Z(w5));   //: @(401,248) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: joint g11 (b) @(332, 176) /w:[ 2 -1 1 4 ]
  //: joint g10 (a) @(301, 154) /w:[ 2 4 1 6 ]
  //: input g6 (b) @(267,176) /sn:0 /w:[ 0 ]
  //: output g9 (Cout) @(560,293) /sn:0 /w:[ 1 ]
  //: input g7 (Cin) @(266,201) /sn:0 /w:[ 0 ]
  //: joint g14 (Cin) @(286, 201) /w:[ 2 -1 1 8 ]
  //: input g5 (a) @(266,154) /sn:0 /w:[ 0 ]
  xor g0 (.I0(a), .I1(b), .I2(Cin), .Z(s));   //: @(407,176) /sn:0 /delay:" 4" /w:[ 3 3 5 0 ]
  //: joint g12 (b) @(332, 295) /w:[ 6 5 -1 8 ]

endmodule

module main;    //: root_module
wire w6;    //: /sn:0 {0}(92,15)(263,15)(263,27){1}
wire w7;    //: /sn:0 {0}(129,347)(129,377)(180,377){1}
wire w16;    //: /sn:0 {0}(92,306)(275,306)(275,326){1}
wire w14;    //: /sn:0 {0}(185,226)(173,226)(173,298)(321,298)(321,378)(311,378){1}
wire w15;    //: /sn:0 {0}(-13,314)(211,314)(211,326){1}
wire w4;    //: /sn:0 {0}(186,-64)(176,-64)(176,9)(320,9)(320,84)(311,84){1}
wire w3;    //: /sn:0 {0}(251,-12)(251,4)(491,4)(491,412)(549,412){1}
wire w0;    //: /sn:0 {0}(-13,-121)(212,-121)(212,-114){1}
wire [3:0] w21;    //: /sn:0 {0}(88,-140)(88,-128){1}
//: {2}(88,-127)(88,14){3}
//: {4}(88,15)(88,155){5}
//: {6}(88,156)(88,305){7}
//: {8}(88,306)(88,516){9}
wire [3:0] w20;    //: /sn:0 {0}(-17,-141)(-17,-122){1}
//: {2}(-17,-121)(-17,20){3}
//: {4}(-17,21)(-17,162){5}
//: {6}(-17,163)(-17,313){7}
//: {8}(-17,314)(-17,502){9}
wire w1;    //: /sn:0 {0}(92,-127)(267,-127)(267,-114){1}
wire w18;    //: /sn:0 /dp:1 {0}(253,442)(253,514)(285,514)(285,448)(383,448)(383,382)(549,382){1}
wire w8;    //: /sn:0 {0}(245,134)(245,145)(478,145)(478,402)(549,402){1}
wire [3:0] w22;    //: /sn:0 /dp:1 {0}(663,340)(663,397)(555,397){1}
wire w12;    //: /sn:0 {0}(373,-100)(383,-100)(383,-60)(311,-60){1}
wire w11;    //: /sn:0 {0}(92,156)(271,156)(271,172){1}
wire w10;    //: /sn:0 {0}(-13,163)(215,163)(215,172){1}
wire w13;    //: /sn:0 /dp:1 {0}(250,286)(250,289)(464,289)(464,392)(549,392){1}
wire w5;    //: /sn:0 {0}(-13,21)(209,21)(209,27){1}
wire w9;    //: /sn:0 {0}(183,79)(173,79)(173,151)(324,151)(324,229)(314,229){1}
//: enddecls

  tran g8(.Z(w15), .I(w20[3]));   //: @(-19,314) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  //: dip g4 (w20) @(-17,-151) /sn:0 /w:[ 0 ] /st:0
  tran g13(.Z(w16), .I(w21[3]));   //: @(86,306) /sn:0 /R:2 /w:[ 0 8 7 ] /ss:1
  FAalterniva g3 (.b(w16), .a(w15), .Cin(w14), .Cout(w7), .s(w18));   //: @(181, 327) /sz:(129, 114) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  FAalterniva g2 (.b(w11), .a(w10), .Cin(w9), .Cout(w14), .s(w13));   //: @(186, 173) /sz:(127, 112) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  FAalterniva g1 (.b(w6), .a(w5), .Cin(w4), .Cout(w9), .s(w8));   //: @(184, 28) /sz:(126, 105) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  led g16 (.I(w7));   //: @(129,340) /sn:0 /w:[ 0 ] /type:0
  tran g11(.Z(w6), .I(w21[1]));   //: @(86,15) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  tran g10(.Z(w1), .I(w21[0]));   //: @(86,-127) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  tran g6(.Z(w5), .I(w20[1]));   //: @(-19,21) /sn:0 /R:2 /w:[ 0 4 3 ] /ss:1
  //: dip g9 (w21) @(88,-150) /sn:0 /w:[ 0 ] /st:0
  tran g7(.Z(w10), .I(w20[2]));   //: @(-19,163) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1
  led g15 (.I(w22));   //: @(663,333) /sn:0 /w:[ 0 ] /type:3
  //: switch g17 (w12) @(356,-100) /sn:0 /w:[ 0 ] /st:0
  concat g14 (.I0(w3), .I1(w8), .I2(w13), .I3(w18), .Z(w22));   //: @(554,397) /sn:0 /w:[ 1 1 1 1 1 ] /dr:0
  tran g5(.Z(w0), .I(w20[0]));   //: @(-19,-121) /sn:0 /R:2 /w:[ 0 2 1 ] /ss:1
  FAalterniva g0 (.b(w1), .a(w0), .Cin(w12), .Cout(w4), .s(w3));   //: @(187, -113) /sz:(123, 100) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  tran g12(.Z(w11), .I(w21[2]));   //: @(86,156) /sn:0 /R:2 /w:[ 0 6 5 ] /ss:1

endmodule

module FAaltern();
//: interface  /sz:(40, 40) /bd:[ ]
//: enddecls


endmodule
