//: version "1.8.7"

module Full_Adder(COut, C, B, A, S);
//: interface  /sz:(40, 40) /bd:[ ]
input B;    //: /sn:0 /dp:1 {0}(240,107)(175,107){1}
//: {2}(171,107)(131,107)(131,151)(96,151){3}
//: {4}(173,109)(173,195)(317,195){5}
input A;    //: /sn:0 {0}(97,102)(142,102){1}
//: {2}(146,102)(240,102){3}
//: {4}(144,104)(144,200)(317,200){5}
output COut;    //: /sn:0 /dp:1 {0}(389,191)(422,191){1}
input C;    //: /sn:0 /dp:1 {0}(345,110)(295,110)(295,176){1}
//: {2}(297,178)(317,178){3}
//: {4}(295,180)(295,198)(95,198){5}
output S;    //: /sn:0 /dp:1 {0}(366,108)(389,108){1}
wire w0;    //: /sn:0 /dp:1 {0}(368,188)(344,188)(344,181)(338,181){1}
wire w1;    //: /sn:0 /dp:1 {0}(368,193)(345,193)(345,198)(338,198){1}
wire w2;    //: /sn:0 {0}(261,105)(274,105){1}
//: {2}(278,105)(345,105){3}
//: {4}(276,107)(276,183)(317,183){5}
//: enddecls

  xor g4 (.I0(w2), .I1(C), .Z(S));   //: @(356,108) /sn:0 /delay:" 4" /w:[ 3 0 0 ]
  and g8 (.I0(B), .I1(A), .Z(w1));   //: @(328,198) /sn:0 /delay:" 3" /w:[ 5 5 1 ]
  //: output g13 (COut) @(419,191) /sn:0 /w:[ 1 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(251,105) /sn:0 /delay:" 4" /w:[ 3 0 0 ]
  //: input g2 (C) @(93,198) /sn:0 /w:[ 5 ]
  //: input g1 (B) @(94,151) /sn:0 /w:[ 3 ]
  or g11 (.I0(w0), .I1(w1), .Z(COut));   //: @(379,191) /sn:0 /delay:" 3" /w:[ 0 0 0 ]
  //: joint g10 (A) @(144, 102) /w:[ 2 -1 1 4 ]
  //: joint g6 (w2) @(276, 105) /w:[ 2 -1 1 4 ]
  //: joint g7 (C) @(295, 178) /w:[ 2 1 -1 4 ]
  //: joint g9 (B) @(173, 107) /w:[ 1 -1 2 4 ]
  and g5 (.I0(C), .I1(w2), .Z(w0));   //: @(328,181) /sn:0 /delay:" 3" /w:[ 3 5 1 ]
  //: input g0 (A) @(95,102) /sn:0 /w:[ 0 ]
  //: output g12 (S) @(386,108) /sn:0 /w:[ 1 ]

endmodule

module CSA(B, S, C, A, COut);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] B;    //: /sn:0 /dp:9 {0}(1,41)(85,41){1}
//: {2}(86,41)(159,41){3}
//: {4}(160,41)(222,41){5}
//: {6}(223,41)(282,41){7}
//: {8}(283,41)(323,41){9}
supply1 w7;    //: /sn:0 /dp:1 {0}(355,160)(370,160){1}
input [3:0] A;    //: /sn:0 /dp:9 {0}(53,25)(103,25){1}
//: {2}(104,25)(176,25){3}
//: {4}(177,25)(246,25){5}
//: {6}(247,25)(305,25){7}
//: {8}(306,25)(315,25){9}
output COut;    //: /sn:0 {0}(-35,157)(-46,157)(-46,118)(-56,118){1}
input C;    //: /sn:0 /dp:3 {0}(-45,318)(18,318){1}
//: {2}(22,318)(154,311)(154,312)(284,312){3}
//: {4}(20,316)(20,117)(-22,117)(-22,134){5}
supply1 w13;    //: /sn:0 {0}(372,98)(318,98){1}
output [3:0] S;    //: /sn:0 {0}(423,336)(307,336)(307,325){1}
wire w6;    //: /sn:0 {0}(215,185)(215,240)(113,240)(113,279){1}
wire S1;    //: /sn:0 {0}(83,180)(83,227)(133,227)(133,279){1}
wire C5;    //: /sn:0 {0}(177,169)(202,169){1}
wire w4;    //: /sn:0 {0}(156,182)(156,233)(123,233)(123,279){1}
wire C6;    //: /sn:0 {0}(109,170)(135,170){1}
wire A3;    //: /sn:0 {0}(104,29)(104,45){1}
//: {2}(102,47)(97,47)(97,66){3}
//: {4}(104,49)(104,138){5}
wire w3;    //: /sn:0 {0}(103,279)(103,247)(285,247)(285,175){1}
wire w0;    //: /sn:0 {0}(306,29)(306,52){1}
//: {2}(308,54)(314,54)(314,133){3}
//: {4}(306,56)(306,65){5}
wire A2;    //: /sn:0 {0}(177,29)(177,47)(169,47){1}
//: {2}(165,47)(161,47)(161,66){3}
//: {4}(167,49)(167,140){5}
wire B2;    //: /sn:0 {0}(160,45)(160,53)(156,53){1}
//: {2}(152,53)(146,53)(146,66){3}
//: {4}(154,55)(154,140){5}
wire C4;    //: /sn:0 {0}(276,168)(244,168){1}
wire w1;    //: /sn:0 {0}(283,45)(283,53){1}
//: {2}(285,55)(294,55)(294,133){3}
//: {4}(283,57)(283,65){5}
wire C2;    //: /sn:0 {0}(177,96)(201,96){1}
wire B1;    //: /sn:0 {0}(223,45)(223,55)(220,55){1}
//: {2}(216,55)(210,55)(210,66){3}
//: {4}(218,57)(218,143){5}
wire w8;    //: /sn:0 /dp:1 {0}(312,250)(312,219)(223,219)(223,108){1}
wire w18;    //: /sn:0 {0}(339,160)(318,160){1}
wire COut2;    //: /sn:0 {0}(135,99)(110,99){1}
wire COut1;    //: /sn:0 {0}(68,98)(4,98)(4,167)(-6,167){1}
wire w11;    //: /sn:0 {0}(332,250)(332,213)(91,213)(91,109){1}
wire w2;    //: /sn:0 {0}(302,107)(302,250){1}
wire w12;    //: /sn:0 {0}(-6,147)(28,147)(28,167)(64,167){1}
wire A1;    //: /sn:0 {0}(247,29)(247,47)(240,47){1}
//: {2}(236,47)(234,47)(234,66){3}
//: {4}(238,49)(238,143){5}
wire B3;    //: /sn:0 {0}(86,45)(86,53){1}
//: {2}(84,55)(77,55)(77,66){3}
//: {4}(86,57)(86,97)(75,97)(75,138){5}
wire C1;    //: /sn:0 {0}(243,98)(274,98){1}
wire [3:0] S3;    //: /sn:0 /dp:1 {0}(118,285)(118,286)(297,286)(297,296){1}
wire [3:0] w9;    //: /sn:0 /dp:1 {0}(317,256)(317,296){1}
wire S2;    //: /sn:0 /dp:1 {0}(162,108)(162,226)(322,226)(322,250){1}
//: enddecls

  concat g4 (.I0(w2), .I1(w8), .I2(S2), .I3(w11), .Z(w9));   //: @(317,255) /sn:0 /R:3 /w:[ 1 0 1 0 0 ] /dr:0
  tran g8(.Z(A2), .I(A[2]));   //: @(177,23) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  tran g13(.Z(B1), .I(B[1]));   //: @(223,39) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  not g37 (.I(w7), .Z(w18));   //: @(349,160) /sn:0 /R:2 /delay:" 4" /w:[ 0 0 ]
  concat g34 (.I0(w3), .I1(w6), .I2(w4), .I3(S1), .Z(S3));   //: @(118,284) /sn:0 /R:3 /w:[ 0 1 1 1 0 ] /dr:0
  Full_Adder g3 (.B(B1), .A(A1), .C(C1), .COut(C2), .S(w8));   //: @(202, 67) /sz:(40, 40) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>0 Lo0<1 Bo0<1 ]
  Full_Adder g2 (.B(w1), .A(w0), .C(w13), .COut(C1), .S(w2));   //: @(275, 66) /sz:(42, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Lo0<1 Bo0<0 ]
  Full_Adder g1 (.B(B2), .A(A2), .C(C2), .COut(COut2), .S(S2));   //: @(136, 67) /sz:(40, 40) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>0 Lo0<0 Bo0<0 ]
  tran g11(.Z(B3), .I(B[3]));   //: @(86,39) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  mux g16 (.I0(S3), .I1(w9), .S(C), .Z(S));   //: @(307,312) /sn:0 /delay:" 2 2" /w:[ 1 1 3 1 ] /ss:0 /do:0
  //: joint g28 (C) @(20, 318) /w:[ 2 4 1 -1 ]
  //: input g10 (B) @(-1,41) /sn:0 /w:[ 0 ]
  //: joint g27 (B2) @(154, 53) /w:[ 1 -1 2 4 ]
  //: output g32 (S) @(420,336) /sn:0 /w:[ 0 ]
  //: input g19 (C) @(-47,318) /sn:0 /w:[ 0 ]
  tran g6(.Z(w0), .I(A[0]));   //: @(306,23) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g7(.Z(A1), .I(A[1]));   //: @(247,23) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g9(.Z(A3), .I(A[3]));   //: @(104,23) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: supply1 g15 (w13) @(372,109) /sn:0 /R:3 /w:[ 0 ]
  //: joint g20 (w1) @(283, 55) /w:[ 2 1 -1 4 ]
  //: joint g31 (A3) @(104, 47) /w:[ -1 1 2 4 ]
  Full_Adder g25 (.B(B2), .A(A2), .C(C5), .COut(C6), .S(w4));   //: @(136, 141) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<1 Bo0<0 ]
  Full_Adder g29 (.B(B3), .A(A3), .C(C6), .COut(w12), .S(S1));   //: @(65, 139) /sz:(43, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<1 Bo0<0 ]
  mux g17 (.I0(w12), .I1(COut1), .S(C), .Z(COut));   //: @(-22,157) /sn:0 /R:3 /delay:" 2 2" /w:[ 0 1 5 0 ] /ss:0 /do:0
  //: input g5 (A) @(51,25) /sn:0 /w:[ 0 ]
  tran g14(.Z(w1), .I(B[0]));   //: @(283,39) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: joint g21 (w0) @(306, 54) /w:[ 2 1 -1 4 ]
  //: supply1 g36 (w7) @(370,171) /sn:0 /R:3 /w:[ 1 ]
  //: joint g24 (A1) @(238, 47) /w:[ 1 -1 2 4 ]
  //: joint g23 (B1) @(218, 55) /w:[ 1 -1 2 4 ]
  Full_Adder g0 (.A(A3), .B(B3), .C(COut2), .COut(COut1), .S(w11));   //: @(69, 67) /sz:(40, 41) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>1 Lo0<0 Bo0<1 ]
  Full_Adder g22 (.A(A1), .B(B1), .C(C4), .COut(C5), .S(w6));   //: @(203, 144) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Lo0<1 Bo0<0 ]
  //: joint g26 (A2) @(167, 47) /w:[ 1 -1 2 4 ]
  tran g12(.Z(B2), .I(B[2]));   //: @(160,39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  Full_Adder g18 (.B(w1), .A(w0), .C(w18), .COut(C4), .S(w3));   //: @(277, 134) /sz:(40, 40) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>1 Lo0<0 Bo0<1 ]
  //: output g33 (COut) @(-53,118) /sn:0 /R:2 /w:[ 1 ]
  //: joint g30 (B3) @(86, 55) /w:[ -1 1 2 4 ]

endmodule

module main;    //: root_module
wire [3:0] B;    //: /sn:0 {0}(113,35)(113,68)(153,68)(153,80){1}
wire [3:0] A;    //: /sn:0 {0}(209,36)(209,69)(167,69)(167,80){1}
wire w0;    //: /sn:0 {0}(97,110)(140,110){1}
wire w1;    //: /sn:0 {0}(182,108)(217,108){1}
wire [3:0] w5;    //: /sn:0 {0}(157,122)(157,163)(180,163){1}
//: enddecls

  led g4 (.I(w1));   //: @(224,108) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: switch g3 (w0) @(80,110) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (A) @(209,26) /sn:0 /w:[ 0 ] /st:13
  //: dip g1 (B) @(113,25) /sn:0 /w:[ 0 ] /st:12
  CSA g6 (.B(B), .A(A), .C(w0), .S(w5), .COut(w1));   //: @(141, 81) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Li0>1 Bo0<0 Ro0<0 ]
  led g5 (.I(w5));   //: @(187,163) /sn:0 /R:3 /w:[ 1 ] /type:3

endmodule
