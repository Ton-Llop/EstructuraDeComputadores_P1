//: version "1.8.7"

module HA(s, b, a, c);
//: interface  /sz:(166, 122) /bd:[ Ti0>a(50/166) Ti1>b(113/166) Lo0<c(59/122) Bo0<s(80/166) ]
input b;    //: /sn:0 {0}(259,188)(281,188){1}
//: {2}(285,188)(321,188)(321,179)(329,179){3}
//: {4}(283,190)(283,235)(330,235){5}
output s;    //: /sn:0 /dp:1 {0}(350,177)(426,177){1}
input a;    //: /sn:0 {0}(260,174)(295,174){1}
//: {2}(299,174)(329,174){3}
//: {4}(297,176)(297,230)(330,230){5}
output c;    //: /sn:0 /dp:1 {0}(351,233)(423,233){1}
//: enddecls

  //: output g4 (s) @(423,177) /sn:0 /w:[ 1 ]
  //: input g3 (b) @(257,188) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(258,174) /sn:0 /w:[ 0 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(341,233) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: joint g6 (a) @(297, 174) /w:[ 2 -1 1 4 ]
  //: joint g7 (b) @(283, 188) /w:[ 2 -1 1 4 ]
  //: output g5 (c) @(420,233) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(340,177) /sn:0 /delay:" 4" /w:[ 3 3 0 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(529,382)(529,387)(498,387)(498,350){1}
wire w0;    //: /sn:0 {0}(469,95)(486,95)(486,156){1}
wire w1;    //: /sn:0 {0}(531,95)(539,95)(539,156){1}
wire w2;    //: /sn:0 {0}(323,231)(323,255)(382,255){1}
wire w5;    //: /sn:0 {0}(401,95)(422,95)(422,156){1}
//: enddecls

  led g4 (.I(w2));   //: @(323,224) /sn:0 /w:[ 0 ] /type:0
  //: switch g3 (w1) @(514,95) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w0) @(452,95) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w5) @(384,95) /sn:0 /w:[ 0 ] /st:0
  led g5 (.I(w4));   //: @(529,375) /sn:0 /w:[ 0 ] /type:0
  FA g0 (.Cin(w1), .b(w0), .a(w5), .Cout(w2), .s(w4));   //: @(383, 157) /sz:(210, 192) /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Lo0<1 Bo0<1 ]

endmodule

module FA(Cin, b, a, Cout, s);
//: interface  /sz:(40, 40) /bd:[ ]
input b;    //: /sn:0 {0}(160,113)(421,113)(421,130){1}
output Cout;    //: /sn:0 /dp:1 {0}(580,442)(700,442){1}
input Cin;    //: /sn:0 {0}(139,250)(582,250)(582,274){1}
output s;    //: /sn:0 /dp:1 {0}(559,378)(559,398)(690,398){1}
input a;    //: /sn:0 {0}(172,96)(382,96)(382,130){1}
wire w0;    //: /sn:0 /dp:1 {0}(559,439)(488,439)(488,324)(505,324){1}
wire w3;    //: /sn:0 {0}(401,230)(401,256)(539,256)(539,274){1}
wire w1;    //: /sn:0 /dp:1 {0}(559,444)(341,444)(341,178)(351,178){1}
//: enddecls

  //: input g4 (Cin) @(137,250) /sn:0 /w:[ 0 ]
  //: input g3 (b) @(158,113) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(170,96) /sn:0 /w:[ 0 ]
  HA g1 (.b(Cin), .a(w3), .c(w0), .s(s));   //: @(506, 275) /sz:(112, 102) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]
  or g6 (.I0(w0), .I1(w1), .Z(Cout));   //: @(570,442) /sn:0 /delay:" 3" /w:[ 0 0 0 ]
  //: output g7 (Cout) @(697,442) /sn:0 /w:[ 1 ]
  //: output g5 (s) @(687,398) /sn:0 /w:[ 1 ]
  HA g0 (.b(b), .a(a), .c(w1), .s(w3));   //: @(352, 131) /sz:(102, 98) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<0 ]

endmodule
