//: version "1.8.7"

module PFA(P, C, B, G, S, A);
//: interface  /sz:(40, 40) /bd:[ ]
input B;    //: /sn:0 {0}(131,81)(169,81){1}
//: {2}(173,81)(240,81)(240,56)(256,56){3}
//: {4}(171,83)(171,175){5}
//: {6}(173,177)(211,177)(211,143)(365,143){7}
//: {8}(171,179)(171,203)(359,203){9}
input A;    //: /sn:0 {0}(134,51)(185,51){1}
//: {2}(189,51)(256,51){3}
//: {4}(187,53)(187,136){5}
//: {6}(189,138)(365,138){7}
//: {8}(187,140)(187,198)(359,198){9}
output G;    //: /sn:0 /dp:1 {0}(380,201)(432,201)(432,190)(487,190){1}
output P;    //: /sn:0 {0}(386,141)(488,141){1}
input C;    //: /sn:0 {0}(121,190)(144,190)(144,153)(247,153)(247,76)(364,76){1}
output S;    //: /sn:0 {0}(385,74)(445,74)(445,97)(482,97){1}
wire w2;    //: /sn:0 {0}(277,54)(314,54)(314,71)(364,71){1}
//: enddecls

  //: output g8 (P) @(485,141) /sn:0 /w:[ 1 ]
  or g4 (.I0(A), .I1(B), .Z(P));   //: @(376,141) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(267,54) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: input g2 (C) @(119,190) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(129,81) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(187, 51) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(w2), .I1(C), .Z(S));   //: @(375,74) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  //: output g9 (G) @(484,190) /sn:0 /w:[ 1 ]
  //: output g7 (S) @(479,97) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(187, 138) /w:[ 6 5 -1 8 ]
  //: joint g11 (B) @(171, 81) /w:[ 2 -1 1 4 ]
  and g5 (.I0(A), .I1(B), .Z(G));   //: @(370,201) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: input g0 (A) @(132,51) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(171, 177) /w:[ 6 5 -1 8 ]

endmodule

module CLA4BITS(C, COut, P, A, B, G, S);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] B;    //: /sn:0 {0}(124,-71)(124,23)(257,23){1}
//: {2}(258,23)(326,23){3}
//: {4}(327,23)(392,23){5}
//: {6}(393,23)(451,23){7}
//: {8}(452,23)(767,23){9}
input [3:0] A;    //: /sn:0 {0}(102,-69)(102,47)(238,47){1}
//: {2}(239,47)(307,47){3}
//: {4}(308,47)(367,47){5}
//: {6}(368,47)(429,47){7}
//: {8}(430,47)(790,47){9}
output G;    //: /sn:0 {0}(432,270)(432,355){1}
output P;    //: /sn:0 {0}(391,270)(391,314)(392,314)(392,341){1}
input C;    //: /sn:0 /dp:3 {0}(466,139)(521,139){1}
//: {2}(525,139)(557,139){3}
//: {4}(523,141)(523,254)(507,254){5}
output COut;    //: /sn:0 {0}(62,251)(176,251)(176,247)(190,247){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(46,186)(94,186){1}
wire w6;    //: /sn:0 {0}(258,27)(258,115){1}
wire w16;    //: /sn:0 /dp:1 {0}(334,155)(334,191)(100,191){1}
wire w13;    //: /sn:0 {0}(341,135)(357,135)(357,228){1}
wire w7;    //: /sn:0 {0}(239,51)(239,59)(241,59)(241,115){1}
wire w4;    //: /sn:0 {0}(308,51)(308,59)(309,59)(309,113){1}
wire w3;    //: /sn:0 {0}(393,27)(393,114){1}
wire w0;    //: /sn:0 {0}(430,51)(430,59)(435,59)(435,116){1}
wire w22;    //: /sn:0 {0}(404,138)(408,138)(408,162)(421,162)(421,207)(430,207)(430,228){1}
wire w20;    //: /sn:0 {0}(460,228)(460,214)(434,214)(434,158){1}
wire w19;    //: /sn:0 {0}(248,157)(248,224)(253,224)(253,228){1}
wire w18;    //: /sn:0 /dp:1 {0}(258,157)(258,201)(100,201){1}
wire w12;    //: /sn:0 {0}(305,155)(305,218)(302,218)(302,228){1}
wire w10;    //: /sn:0 {0}(458,158)(458,171)(100,171){1}
wire w23;    //: /sn:0 {0}(270,134)(287,134)(287,228){1}
wire w21;    //: /sn:0 {0}(487,228)(487,217)(463,217)(463,187)(445,187)(445,158){1}
wire w1;    //: /sn:0 {0}(452,27)(452,35)(455,35)(455,116){1}
wire w8;    //: /sn:0 {0}(367,228)(367,215)(370,215)(370,156){1}
wire w14;    //: /sn:0 {0}(394,156)(394,181)(100,181){1}
wire w2;    //: /sn:0 {0}(368,51)(368,59)(371,59)(371,114){1}
wire w11;    //: /sn:0 {0}(226,228)(226,180)(236,180)(236,157){1}
wire w15;    //: /sn:0 {0}(321,155)(321,228){1}
wire w5;    //: /sn:0 {0}(327,27)(327,35)(328,35)(328,113){1}
wire w9;    //: /sn:0 {0}(389,228)(389,200)(381,200)(381,156){1}
//: enddecls

  //: input g4 (C) @(559,139) /sn:0 /R:2 /w:[ 3 ]
  tran g8(.Z(w7), .I(A[3]));   //: @(239,45) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  PFA g3 (.B(w1), .A(w0), .C(C), .S(w10), .G(w21), .P(w20));   //: @(425, 117) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<1 ]
  //: joint g16 (C) @(523, 139) /w:[ 2 -1 1 4 ]
  //: output g17 (COut) @(65,251) /sn:0 /R:2 /w:[ 0 ]
  PFA g2 (.B(w3), .A(w2), .C(w22), .S(w14), .G(w9), .P(w8));   //: @(363, 115) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<1 ]
  PFA g1 (.B(w5), .A(w4), .C(w13), .S(w16), .G(w15), .P(w12));   //: @(300, 114) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g18 (P) @(392,338) /sn:0 /R:3 /w:[ 1 ]
  tran g10(.Z(w4), .I(A[2]));   //: @(308,45) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: input g6 (A) @(102,-71) /sn:0 /R:3 /w:[ 0 ]
  //: input g7 (B) @(124,-73) /sn:0 /R:3 /w:[ 0 ]
  tran g9(.Z(w6), .I(B[3]));   //: @(258,21) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g12(.Z(w2), .I(A[1]));   //: @(368,45) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g11(.Z(w5), .I(B[2]));   //: @(327,21) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  CLALogic g5 (.G3(w19), .P3(w11), .G2(w15), .P2(w12), .G1(w9), .P1(w8), .G0(w21), .P0(w20), .C0(C), .C3(w23), .C1(w22), .C2(w13), .C4(COut), .GG(G), .PG(P));   //: @(191, 229) /sz:(315, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>1 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 To0<1 To1<1 To2<1 Lo0<1 Bo0<0 Bo1<0 ]
  tran g14(.Z(w0), .I(A[0]));   //: @(430,45) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: output g19 (G) @(432,352) /sn:0 /R:3 /w:[ 1 ]
  //: output g21 (S) @(49,186) /sn:0 /R:2 /w:[ 0 ]
  concat g20 (.I0(w10), .I1(w14), .I2(w16), .I3(w18), .Z(S));   //: @(95,186) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0
  tran g15(.Z(w1), .I(B[0]));   //: @(452,21) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  PFA g0 (.B(w6), .A(w7), .C(w23), .S(w18), .G(w19), .P(w11));   //: @(229, 116) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<0 Bo2<1 ]
  tran g13(.Z(w3), .I(B[1]));   //: @(393,21) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1

endmodule

module CLALogic(G2, C4, P2, P0, G3, G0, C3, P1, G1, P3, GG, C1, C2, C0, PG);
//: interface  /sz:(40, 40) /bd:[ ]
input G2;    //: /sn:0 {0}(138,533)(192,533){1}
//: {2}(196,533)(410,533){3}
//: {4}(414,533)(739,533)(739,445)(747,445){5}
//: {6}(412,535)(412,580)(491,580){7}
//: {8}(194,535)(194,908)(639,908){9}
input C0;    //: /sn:0 /dp:3 {0}(381,117)(332,117){1}
//: {2}(328,117)(237,117){3}
//: {4}(233,117)(181,117){5}
//: {6}(177,117)(148,117)(148,139)(144,139){7}
//: {8}(179,119)(179,748)(496,748){9}
//: {10}(235,119)(235,474)(563,474){11}
//: {12}(330,119)(330,220)(407,220){13}
output GG;    //: /sn:0 /dp:1 {0}(841,936)(934,936)(934,937)(946,937){1}
input P1;    //: /sn:0 {0}(654,864)(305,864)(305,271){1}
//: {2}(307,269)(386,269)(386,263)(392,263){3}
//: {4}(303,269)(292,269){5}
//: {6}(288,269)(262,269){7}
//: {8}(258,269)(247,269){9}
//: {10}(243,269)(209,269){11}
//: {12}(205,269)(177,269){13}
//: {14}(175,267)(175,263)(153,263)(153,301)(198,301)(198,429)(552,429){15}
//: {16}(173,269)(142,269){17}
//: {18}(175,271)(175,484)(563,484){19}
//: {20}(207,271)(207,713)(496,713){21}
//: {22}(245,271)(245,753)(496,753){23}
//: {24}(260,271)(260,281)(268,281)(268,989)(649,989){25}
//: {26}(290,271)(290,339)(320,339)(320,230)(407,230){27}
output C3;    //: /sn:0 /dp:1 {0}(903,445)(849,445)(849,437)(768,437){1}
output PG;    //: /sn:0 {0}(675,861)(936,861){1}
input G0;    //: /sn:0 /dp:9 {0}(141,170)(216,170){1}
//: {2}(220,170)(250,170){3}
//: {4}(254,170)(270,170){5}
//: {6}(274,170)(301,170){7}
//: {8}(305,170)(648,170)(648,148)(600,148)(600,133)(606,133){9}
//: {10}(303,172)(303,984)(649,984){11}
//: {12}(272,172)(272,258)(392,258){13}
//: {14}(252,172)(252,703)(496,703){15}
//: {16}(218,172)(218,424)(552,424){17}
output C4;    //: /sn:0 {0}(708,694)(927,694){1}
output C2;    //: /sn:0 {0}(623,261)(770,261)(770,262)(780,262){1}
input P3;    //: /sn:0 {0}(643,951)(206,951)(206,740){1}
//: {2}(208,738)(260,738)(260,763)(496,763){3}
//: {4}(204,738)(167,738){5}
//: {6}(165,736)(165,585)(491,585){7}
//: {8}(163,738)(151,738){9}
//: {10}(147,738)(126,738){11}
//: {12}(124,736)(124,718)(496,718){13}
//: {14}(122,738)(108,738){15}
//: {16}(106,736)(106,726)(121,726)(121,999)(649,999){17}
//: {18}(104,738)(93,738){19}
//: {20}(106,740)(106,869)(654,869){21}
//: {22}(124,740)(124,750)(139,750)(139,659)(499,659){23}
//: {24}(149,740)(149,903)(639,903){25}
input G1;    //: /sn:0 /dp:11 {0}(148,311)(271,311){1}
//: {2}(275,311)(370,311){3}
//: {4}(374,311)(455,311){5}
//: {6}(459,311)(594,311)(594,266)(602,266){7}
//: {8}(457,313)(457,381)(557,381){9}
//: {10}(372,313)(372,941)(643,941){11}
//: {12}(273,313)(273,649)(499,649){13}
input G3;    //: /sn:0 {0}(89,801)(250,801){1}
//: {2}(254,801)(645,801)(645,704)(687,704){3}
//: {4}(252,803)(252,934)(820,934){5}
output C1;    //: /sn:0 {0}(627,131)(770,131){1}
input P0;    //: /sn:0 {0}(145,106)(195,106){1}
//: {2}(199,106)(217,106){3}
//: {4}(221,106)(286,106){5}
//: {6}(290,106)(344,106){7}
//: {8}(348,106)(377,106)(377,112)(381,112){9}
//: {10}(346,108)(346,854)(654,854){11}
//: {12}(288,108)(288,225)(407,225){13}
//: {14}(219,108)(219,743)(496,743){15}
//: {16}(197,108)(197,479)(563,479){17}
input P2;    //: /sn:0 /dp:21 {0}(649,994)(182,994)(182,432){1}
//: {2}(184,430)(212,430){3}
//: {4}(216,430)(294,430){5}
//: {6}(298,430)(356,430)(356,489)(563,489){7}
//: {8}(296,432)(296,466)(310,466)(310,434)(552,434){9}
//: {10}(214,428)(214,386)(557,386){11}
//: {12}(180,430)(158,430){13}
//: {14}(156,428)(156,418)(171,418)(171,708)(496,708){15}
//: {16}(154,430)(142,430){17}
//: {18}(140,428)(140,377)(160,377)(160,391)(171,391)(171,416)(187,416){19}
//: {20}(191,416)(293,416)(293,859)(654,859){21}
//: {22}(189,418)(189,946)(643,946){23}
//: {24}(138,430)(127,430){25}
//: {26}(140,432)(140,654)(499,654){27}
//: {28}(156,432)(156,758)(496,758){29}
wire w6;    //: /sn:0 {0}(578,384)(737,384)(737,430)(747,430){1}
wire w16;    //: /sn:0 {0}(820,939)(674,939)(674,946)(664,946){1}
wire w7;    //: /sn:0 {0}(413,261)(602,261){1}
wire w4;    //: /sn:0 {0}(517,753)(634,753)(634,699)(687,699){1}
wire w0;    //: /sn:0 /dp:1 {0}(820,929)(670,929)(670,906)(660,906){1}
wire w3;    //: /sn:0 {0}(428,225)(592,225)(592,256)(602,256){1}
wire w12;    //: /sn:0 {0}(512,583)(677,583)(677,684)(687,684){1}
wire w10;    //: /sn:0 {0}(517,710)(584,710)(584,694)(687,694){1}
wire w17;    //: /sn:0 {0}(820,944)(680,944)(680,991)(670,991){1}
wire w2;    //: /sn:0 {0}(402,115)(596,115)(596,128)(606,128){1}
wire w11;    //: /sn:0 {0}(520,654)(593,654)(593,681)(656,681)(656,689)(687,689){1}
wire w5;    //: /sn:0 {0}(573,429)(719,429)(719,435)(747,435){1}
wire w9;    //: /sn:0 {0}(747,440)(594,440)(594,481)(584,481){1}
//: enddecls

  or g4 (.I0(w2), .I1(G0), .Z(C1));   //: @(617,131) /sn:0 /delay:" 3" /w:[ 1 9 0 ]
  and g8 (.I0(C0), .I1(P0), .I2(P1), .Z(w3));   //: @(418,225) /sn:0 /delay:" 3" /w:[ 13 13 27 0 ]
  //: joint g44 (P3) @(165, 738) /w:[ 5 6 8 -1 ]
  and g3 (.I0(P0), .I1(C0), .Z(w2));   //: @(392,115) /sn:0 /delay:" 3" /w:[ 9 0 0 ]
  //: input g16 (G2) @(136,533) /sn:0 /w:[ 0 ]
  //: output g47 (C4) @(924,694) /sn:0 /w:[ 1 ]
  //: input g17 (P2) @(125,430) /sn:0 /w:[ 25 ]
  //: joint g26 (G1) @(457, 311) /w:[ 6 -1 5 8 ]
  //: input g2 (P0) @(143,106) /sn:0 /w:[ 0 ]
  //: joint g23 (G0) @(218, 170) /w:[ 2 -1 1 16 ]
  //: input g30 (G3) @(87,801) /sn:0 /w:[ 0 ]
  //: input g1 (G0) @(139,170) /sn:0 /w:[ 0 ]
  //: joint g39 (P3) @(124, 738) /w:[ 11 12 14 22 ]
  //: joint g24 (P2) @(296, 430) /w:[ 6 -1 5 8 ]
  //: output g29 (C3) @(900,445) /sn:0 /w:[ 0 ]
  //: joint g60 (G1) @(372, 311) /w:[ 4 -1 3 10 ]
  //: joint g51 (P1) @(305, 269) /w:[ 2 -1 4 1 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w9));   //: @(574,481) /sn:0 /delay:" 3" /w:[ 11 17 19 7 1 ]
  or g65 (.I0(w0), .I1(G3), .I2(w16), .I3(w17), .Z(GG));   //: @(831,936) /sn:0 /delay:" 3" /w:[ 0 5 0 0 0 ]
  //: joint g10 (G0) @(272, 170) /w:[ 6 -1 5 12 ]
  and g25 (.I0(G1), .I1(P2), .Z(w6));   //: @(568,384) /sn:0 /delay:" 3" /w:[ 9 11 0 ]
  //: joint g64 (G0) @(303, 170) /w:[ 8 -1 7 10 ]
  and g49 (.I0(P0), .I1(P2), .I2(P1), .I3(P3), .Z(PG));   //: @(665,861) /sn:0 /delay:" 3" /w:[ 11 21 0 21 0 ]
  //: joint g50 (P0) @(346, 106) /w:[ 8 -1 7 10 ]
  //: input g6 (P1) @(140,269) /sn:0 /w:[ 17 ]
  //: joint g58 (P3) @(206, 738) /w:[ 2 -1 4 1 ]
  //: input g7 (G1) @(146,311) /sn:0 /w:[ 0 ]
  and g9 (.I0(G0), .I1(P1), .Z(w7));   //: @(403,261) /sn:0 /delay:" 3" /w:[ 13 3 0 ]
  //: joint g56 (G2) @(194, 533) /w:[ 2 -1 1 8 ]
  //: joint g35 (P2) @(156, 430) /w:[ 13 14 16 28 ]
  //: joint g59 (P2) @(189, 416) /w:[ 20 -1 19 22 ]
  //: input g31 (P3) @(91,738) /sn:0 /w:[ 19 ]
  and g22 (.I0(G0), .I1(P1), .I2(P2), .Z(w5));   //: @(563,429) /sn:0 /delay:" 3" /w:[ 17 15 9 0 ]
  //: output g67 (GG) @(943,937) /sn:0 /w:[ 1 ]
  and g36 (.I0(G0), .I1(P2), .I2(P1), .I3(P3), .Z(w10));   //: @(507,710) /sn:0 /delay:" 3" /w:[ 15 15 21 13 0 ]
  //: joint g41 (G1) @(273, 311) /w:[ 2 -1 1 12 ]
  and g54 (.I0(P3), .I1(G2), .Z(w0));   //: @(650,906) /sn:0 /delay:" 3" /w:[ 25 9 1 ]
  //: joint g45 (G2) @(412, 533) /w:[ 4 -1 3 6 ]
  //: joint g33 (P0) @(219, 106) /w:[ 4 -1 3 14 ]
  //: joint g42 (P2) @(140, 430) /w:[ 17 18 24 26 ]
  //: joint g52 (P3) @(106, 738) /w:[ 15 16 18 20 ]
  and g40 (.I0(G1), .I1(P2), .I2(P3), .Z(w11));   //: @(510,654) /sn:0 /delay:" 3" /w:[ 13 27 23 0 ]
  //: joint g66 (G3) @(252, 801) /w:[ 2 -1 1 4 ]
  //: joint g12 (C0) @(330, 117) /w:[ 1 -1 2 12 ]
  //: joint g34 (P1) @(245, 269) /w:[ 9 -1 10 22 ]
  or g28 (.I0(w6), .I1(w5), .I2(w9), .I3(G2), .Z(C3));   //: @(758,437) /sn:0 /delay:" 3" /w:[ 1 1 0 5 1 ]
  and g57 (.I0(G1), .I1(P2), .I2(P3), .Z(w16));   //: @(654,946) /sn:0 /delay:" 3" /w:[ 11 23 0 1 ]
  or g46 (.I0(w12), .I1(w11), .I2(w10), .I3(w4), .I4(G3), .Z(C4));   //: @(698,694) /sn:0 /delay:" 3" /w:[ 1 1 1 1 3 0 ]
  //: joint g11 (P0) @(288, 106) /w:[ 6 -1 5 12 ]
  //: output g5 (C1) @(767,131) /sn:0 /w:[ 1 ]
  or g14 (.I0(w3), .I1(w7), .I2(G1), .Z(C2));   //: @(613,261) /sn:0 /delay:" 3" /w:[ 1 1 7 0 ]
  and g61 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w17));   //: @(660,991) /sn:0 /delay:" 3" /w:[ 11 25 0 17 1 ]
  //: joint g19 (C0) @(235, 117) /w:[ 3 -1 4 10 ]
  //: joint g21 (P1) @(175, 269) /w:[ 13 14 16 18 ]
  and g32 (.I0(P0), .I1(C0), .I2(P1), .I3(P2), .I4(P3), .Z(w4));   //: @(507,753) /sn:0 /delay:" 3" /w:[ 15 9 23 29 3 0 ]
  //: joint g20 (P0) @(197, 106) /w:[ 2 -1 1 16 ]
  //: joint g63 (P1) @(260, 269) /w:[ 7 -1 8 24 ]
  //: joint g38 (P1) @(207, 269) /w:[ 11 -1 12 20 ]
  //: output g15 (C2) @(777,262) /sn:0 /w:[ 1 ]
  and g43 (.I0(G2), .I1(P3), .Z(w12));   //: @(502,583) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: input g0 (C0) @(142,139) /sn:0 /w:[ 7 ]
  //: joint g27 (P2) @(214, 430) /w:[ 4 10 3 -1 ]
  //: joint g48 (C0) @(179, 117) /w:[ 5 -1 6 8 ]
  //: joint g37 (G0) @(252, 170) /w:[ 4 -1 3 14 ]
  //: joint g62 (P2) @(182, 430) /w:[ 2 -1 12 1 ]
  //: joint g55 (P3) @(149, 738) /w:[ 9 -1 10 24 ]
  //: joint g13 (P1) @(290, 269) /w:[ 5 -1 6 26 ]
  //: output g53 (PG) @(933,861) /sn:0 /w:[ 1 ]

endmodule

module main;    //: root_module
wire w7;    //: /sn:0 {0}(256,305)(336,305)(336,293)(399,293){1}
wire [3:0] w4;    //: /sn:0 {0}(378,97)(378,139)(416,139)(416,146)(433,146)(433,203){1}
wire [3:0] w0;    //: /sn:0 {0}(481,336)(481,469)(593,469)(593,459){1}
wire [3:0] w3;    //: /sn:0 /dp:1 {0}(519,203)(519,147)(535,147)(535,84){1}
wire w1;    //: /sn:0 /dp:1 {0}(564,268)(744,268){1}
wire w8;    //: /sn:0 {0}(249,221)(389,221)(389,231)(399,231){1}
wire w5;    //: /sn:0 {0}(249,269)(276,269)(276,270)(399,270){1}
//: enddecls

  //: dip g4 (w4) @(378,87) /sn:0 /w:[ 0 ] /st:15
  led g3 (.I(w5));   //: @(242,269) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: switch g2 (w1) @(762,268) /sn:0 /R:2 /w:[ 1 ] /st:0
  led g1 (.I(w0));   //: @(593,452) /sn:0 /w:[ 1 ] /type:3
  led g6 (.I(w7));   //: @(249,305) /sn:0 /R:1 /w:[ 0 ] /type:0
  led g7 (.I(w8));   //: @(242,221) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: dip g5 (w3) @(535,74) /sn:0 /w:[ 1 ] /st:15
  CLA4BITS g0 (.B(w3), .A(w4), .C(w1), .G(w8), .P(w7), .COut(w5), .S(w0));   //: @(400, 204) /sz:(163, 131) /sn:0 /p:[ Ti0>0 Ti1>1 Ri0>0 Lo0<1 Lo1<1 Lo2<1 Bo0<0 ]

endmodule
