//: version "1.8.7"

module CLA16BITS(C, COut, P, A, B, S, G);
//: interface  /sz:(40, 40) /bd:[ ]
input [15:0] B;    //: /sn:0 {0}(144,-51)(144,43)(277,43){1}
//: {2}(278,43)(346,43){3}
//: {4}(347,43)(412,43){5}
//: {6}(413,43)(471,43){7}
//: {8}(472,43)(787,43){9}
input [15:0] A;    //: /sn:0 {0}(122,-49)(122,67)(258,67){1}
//: {2}(259,67)(327,67){3}
//: {4}(328,67)(387,67){5}
//: {6}(388,67)(449,67){7}
//: {8}(450,67)(810,67){9}
output G;    //: /sn:0 {0}(446,434)(446,348){1}
output P;    //: /sn:0 {0}(396,348)(396,393)(395,393)(395,439){1}
input C;    //: /sn:0 {0}(574,139)(558,139)(558,145)(536,145){1}
//: {2}(532,145)(506,145)(506,143)(482,143){3}
//: {4}(534,147)(534,322)(507,322){5}
output COut;    //: /sn:0 /dp:1 {0}(82,271)(182,271)(182,324)(206,324){1}
output [15:0] S;    //: /sn:0 {0}(66,206)(114,206){1}
wire w13;    //: /sn:0 /dp:1 {0}(265,288)(265,275)(267,275)(267,163){1}
wire [3:0] w6;    //: /sn:0 {0}(278,47)(278,111)(273,111)(273,121){1}
wire [3:0] w7;    //: /sn:0 {0}(259,71)(259,111)(258,111)(258,121){1}
wire [3:0] w4;    //: /sn:0 {0}(328,71)(328,82)(322,82)(322,113){1}
wire [3:0] w36;    //: /sn:0 {0}(342,155)(342,172)(349,172)(349,211)(120,211){1}
wire [3:0] w0;    //: /sn:0 {0}(450,71)(450,109)(454,109)(454,119){1}
wire [3:0] w3;    //: /sn:0 {0}(413,47)(413,110)(408,110)(408,120){1}
wire w20;    //: /sn:0 {0}(448,162)(448,239)(471,239)(471,288){1}
wire w12;    //: /sn:0 /dp:1 {0}(316,155)(316,284)(315,284)(315,288){1}
wire [3:0] w10;    //: /sn:0 {0}(120,191)(474,191)(474,162){1}
wire w23;    //: /sn:0 /dp:1 {0}(289,142)(309,142)(309,150)(298,150)(298,288){1}
wire w21;    //: /sn:0 {0}(462,162)(462,212)(454,212)(454,242)(480,242)(480,288){1}
wire [3:0] w1;    //: /sn:0 {0}(472,47)(472,109)(471,109)(471,119){1}
wire w31;    //: /sn:0 /dp:1 {0}(251,163)(251,256)(236,256)(236,288){1}
wire w8;    //: /sn:0 {0}(350,133)(369,133)(369,288){1}
wire [3:0] w46;    //: /sn:0 {0}(414,162)(414,201)(120,201){1}
wire [3:0] w33;    //: /sn:0 {0}(280,163)(280,221)(120,221){1}
wire w48;    //: /sn:0 /dp:1 {0}(388,162)(388,265)(393,265)(393,288){1}
wire w11;    //: /sn:0 {0}(333,288)(333,212)(330,212)(330,155){1}
wire [3:0] w2;    //: /sn:0 {0}(388,71)(388,112)(394,112)(394,120){1}
wire w47;    //: /sn:0 /dp:1 {0}(402,162)(402,250)(414,250)(414,288){1}
wire [3:0] w5;    //: /sn:0 {0}(347,47)(347,109)(336,109)(336,113){1}
wire w9;    //: /sn:0 {0}(422,140)(434,140)(434,164)(422,164)(422,228)(448,228)(448,288){1}
//: enddecls

  //: input g4 (C) @(576,139) /sn:0 /R:2 /w:[ 0 ]
  tran g8(.Z(w7), .I(A[15:12]));   //: @(259,65) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: output g17 (COut) @(85,271) /sn:0 /R:2 /w:[ 0 ]
  //: joint g2 (C) @(534, 145) /w:[ 1 -1 2 4 ]
  CLA4BITS g23 (.B(w1), .A(w0), .C(C), .S(w10), .G(w21), .P(w20));   //: @(441, 120) /sz:(40, 41) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>3 Bo0<1 Bo1<0 Bo2<0 ]
  CLA4BITS g24 (.B(w3), .A(w2), .C(w9), .S(w46), .G(w47), .P(w48));   //: @(381, 121) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<0 Bo2<0 ]
  CLA4BITS g1 (.B(w6), .A(w7), .C(w23), .S(w33), .G(w13), .P(w31));   //: @(244, 122) /sz:(44, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<0 ]
  //: output g18 (P) @(395,436) /sn:0 /R:3 /w:[ 1 ]
  tran g10(.Z(w4), .I(A[11:8]));   //: @(328,65) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: input g6 (A) @(122,-51) /sn:0 /R:3 /w:[ 0 ]
  //: input g7 (B) @(144,-53) /sn:0 /R:3 /w:[ 0 ]
  tran g9(.Z(w6), .I(B[15:12]));   //: @(278,41) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  CLA4BITS g22 (.B(w5), .A(w4), .C(w8), .S(w36), .G(w11), .P(w12));   //: @(309, 114) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<0 ]
  tran g12(.Z(w2), .I(A[7:4]));   //: @(388,65) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  tran g14(.Z(w0), .I(A[3:0]));   //: @(450,65) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g11(.Z(w5), .I(B[11:8]));   //: @(347,41) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: output g21 (S) @(69,206) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (G) @(446,431) /sn:0 /R:3 /w:[ 0 ]
  concat g20 (.I0(w10), .I1(w46), .I2(w36), .I3(w33), .Z(S));   //: @(115,206) /sn:0 /R:2 /w:[ 0 1 1 1 1 ] /dr:0
  LookaheadCarryUnit g0 (.G8(w11), .P12(w31), .G12(w13), .P8(w12), .G4(w47), .P4(w48), .G0(w21), .P0(w20), .C0(C), .C8(w8), .C12(w23), .C4(w9), .C16(COut), .GG(G), .PG(P));   //: @(207, 289) /sz:(299, 58) /sn:0 /p:[ Ti0>0 Ti1>1 Ti2>0 Ti3>1 Ti4>1 Ti5>1 Ti6>1 Ti7>1 Ri0>5 To0<1 To1<1 To2<1 Lo0<1 Bo0<1 Bo1<0 ]
  tran g15(.Z(w1), .I(B[3:0]));   //: @(472,41) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g13(.Z(w3), .I(B[7:4]));   //: @(413,41) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1

endmodule

module PFA(P, C, B, G, S, A);
//: interface  /sz:(40, 40) /bd:[ ]
input B;    //: /sn:0 {0}(131,81)(169,81){1}
//: {2}(173,81)(236,81)(236,56)(252,56){3}
//: {4}(171,83)(171,175){5}
//: {6}(173,177)(216,177)(216,143)(370,143){7}
//: {8}(171,179)(171,203)(359,203){9}
input A;    //: /sn:0 {0}(134,51)(185,51){1}
//: {2}(189,51)(252,51){3}
//: {4}(187,53)(187,136){5}
//: {6}(189,138)(370,138){7}
//: {8}(187,140)(187,198)(359,198){9}
output G;    //: /sn:0 /dp:1 {0}(380,201)(432,201)(432,190)(487,190){1}
output P;    //: /sn:0 {0}(391,141)(488,141){1}
input C;    //: /sn:0 {0}(121,190)(144,190)(144,153)(247,153)(247,76)(364,76){1}
output S;    //: /sn:0 {0}(385,74)(445,74)(445,97)(482,97){1}
wire w2;    //: /sn:0 {0}(273,54)(310,54)(310,71)(364,71){1}
//: enddecls

  //: output g8 (P) @(485,141) /sn:0 /w:[ 1 ]
  or g4 (.I0(A), .I1(B), .Z(P));   //: @(381,141) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(263,54) /sn:0 /delay:" 4" /w:[ 3 3 0 ]
  //: input g2 (C) @(119,190) /sn:0 /w:[ 0 ]
  //: input g1 (B) @(129,81) /sn:0 /w:[ 0 ]
  //: joint g10 (A) @(187, 51) /w:[ 2 -1 1 4 ]
  xor g6 (.I0(w2), .I1(C), .Z(S));   //: @(375,74) /sn:0 /delay:" 4" /w:[ 1 1 0 ]
  //: output g9 (G) @(484,190) /sn:0 /w:[ 1 ]
  //: output g7 (S) @(479,97) /sn:0 /w:[ 1 ]
  //: joint g12 (A) @(187, 138) /w:[ 6 5 -1 8 ]
  and g5 (.I0(A), .I1(B), .Z(G));   //: @(370,201) /sn:0 /delay:" 3" /w:[ 9 9 0 ]
  //: joint g11 (B) @(171, 81) /w:[ 2 -1 1 4 ]
  //: input g0 (A) @(132,51) /sn:0 /w:[ 0 ]
  //: joint g13 (B) @(171, 177) /w:[ 6 5 -1 8 ]

endmodule

module LookaheadCarryUnit(C16, G8, P8, P0, G12, G0, C12, P4, G4, P12, GG, C4, C0, C8, PG);
//: interface  /sz:(40, 40) /bd:[ ]
input P4;    //: /sn:0 /dp:26 {0}(673,884)(324,884)(324,291){1}
//: {2}(326,289)(405,289)(405,283)(411,283){3}
//: {4}(322,289)(311,289){5}
//: {6}(307,289)(281,289){7}
//: {8}(277,289)(266,289){9}
//: {10}(262,289)(228,289){11}
//: {12}(224,289)(196,289){13}
//: {14}(194,287)(194,283)(172,283)(172,321)(217,321)(217,449)(571,449){15}
//: {16}(192,289)(161,289){17}
//: {18}(194,291)(194,504)(582,504){19}
//: {20}(226,291)(226,733)(515,733){21}
//: {22}(264,291)(264,773)(515,773){23}
//: {24}(279,291)(279,301)(288,301)(288,1009)(670,1009){25}
//: {26}(309,291)(309,359)(339,359)(339,250)(426,250){27}
output C12;    //: /sn:0 {0}(922,465)(868,465)(868,457)(787,457){1}
input P8;    //: /sn:0 /dp:25 {0}(670,1014)(201,1014)(201,452){1}
//: {2}(203,450)(231,450){3}
//: {4}(235,450)(313,450){5}
//: {6}(317,450)(375,450)(375,509)(582,509){7}
//: {8}(315,452)(315,486)(329,486)(329,454)(571,454){9}
//: {10}(233,448)(233,406)(576,406){11}
//: {12}(199,450)(177,450){13}
//: {14}(175,448)(175,438)(190,438)(190,728)(515,728){15}
//: {16}(173,450)(161,450){17}
//: {18}(159,448)(159,397)(179,397)(179,411)(190,411)(190,436)(206,436){19}
//: {20}(210,436)(312,436)(312,879)(673,879){21}
//: {22}(208,438)(208,966)(662,966){23}
//: {24}(157,450)(146,450){25}
//: {26}(159,452)(159,674)(518,674){27}
//: {28}(175,452)(175,778)(515,778){29}
output GG;    //: /sn:0 {0}(861,956)(954,956)(954,957)(966,957){1}
input C0;    //: /sn:0 {0}(400,137)(351,137){1}
//: {2}(347,137)(256,137){3}
//: {4}(252,137)(200,137){5}
//: {6}(196,137)(167,137)(167,159)(163,159){7}
//: {8}(198,139)(198,768)(515,768){9}
//: {10}(254,139)(254,494)(582,494){11}
//: {12}(349,139)(349,240)(426,240){13}
input G8;    //: /sn:0 {0}(135,550)(162,550)(162,553)(211,553){1}
//: {2}(215,553)(429,553){3}
//: {4}(433,553)(758,553)(758,465)(766,465){5}
//: {6}(431,555)(431,600)(510,600){7}
//: {8}(213,555)(213,928)(658,928){9}
output C16;    //: /sn:0 /dp:1 {0}(727,714)(946,714){1}
output PG;    //: /sn:0 {0}(694,881)(956,881){1}
input G0;    //: /sn:0 {0}(160,190)(235,190){1}
//: {2}(239,190)(269,190){3}
//: {4}(273,190)(289,190){5}
//: {6}(293,190)(320,190){7}
//: {8}(324,190)(667,190)(667,168)(619,168)(619,153)(625,153){9}
//: {10}(322,192)(322,1004)(670,1004){11}
//: {12}(291,192)(291,278)(411,278){13}
//: {14}(271,192)(271,723)(515,723){15}
//: {16}(237,192)(237,444)(571,444){17}
output C4;    //: /sn:0 /dp:1 {0}(646,151)(789,151){1}
input G4;    //: /sn:0 {0}(167,331)(290,331){1}
//: {2}(294,331)(389,331){3}
//: {4}(393,331)(474,331){5}
//: {6}(478,331)(613,331)(613,286)(621,286){7}
//: {8}(476,333)(476,401)(576,401){9}
//: {10}(391,333)(391,961)(662,961){11}
//: {12}(292,333)(292,669)(518,669){13}
input P12;    //: /sn:0 {0}(662,971)(225,971)(225,760){1}
//: {2}(227,758)(279,758)(279,783)(515,783){3}
//: {4}(223,758)(186,758){5}
//: {6}(184,756)(184,605)(510,605){7}
//: {8}(182,758)(170,758){9}
//: {10}(166,758)(145,758){11}
//: {12}(143,756)(143,738)(515,738){13}
//: {14}(141,758)(127,758){15}
//: {16}(125,756)(125,746)(141,746)(141,1019)(670,1019){17}
//: {18}(123,758)(112,758){19}
//: {20}(125,760)(125,889)(673,889){21}
//: {22}(143,760)(143,770)(158,770)(158,679)(518,679){23}
//: {24}(168,760)(168,923)(658,923){25}
input P0;    //: /sn:0 {0}(164,126)(214,126){1}
//: {2}(218,126)(236,126){3}
//: {4}(240,126)(305,126){5}
//: {6}(309,126)(363,126){7}
//: {8}(367,126)(394,126)(394,132)(400,132){9}
//: {10}(365,128)(365,874)(673,874){11}
//: {12}(307,128)(307,245)(426,245){13}
//: {14}(238,128)(238,763)(515,763){15}
//: {16}(216,128)(216,499)(582,499){17}
output C8;    //: /sn:0 /dp:1 {0}(642,281)(789,281)(789,282)(799,282){1}
input G12;    //: /sn:0 {0}(108,821)(258,821){1}
//: {2}(262,821)(664,821)(664,724)(706,724){3}
//: {4}(260,823)(260,954)(840,954){5}
wire w16;    //: /sn:0 {0}(840,959)(693,959)(693,966)(683,966){1}
wire w6;    //: /sn:0 {0}(597,404)(756,404)(756,450)(766,450){1}
wire w7;    //: /sn:0 {0}(432,281)(621,281){1}
wire w4;    //: /sn:0 {0}(536,773)(653,773)(653,719)(706,719){1}
wire w0;    //: /sn:0 {0}(840,949)(689,949)(689,926)(679,926){1}
wire w3;    //: /sn:0 {0}(447,245)(611,245)(611,276)(621,276){1}
wire w12;    //: /sn:0 {0}(531,603)(696,603)(696,704)(706,704){1}
wire w10;    //: /sn:0 {0}(536,730)(603,730)(603,714)(706,714){1}
wire w17;    //: /sn:0 {0}(840,964)(701,964)(701,1011)(691,1011){1}
wire w11;    //: /sn:0 /dp:1 {0}(539,674)(612,674)(612,701)(675,701)(675,709)(706,709){1}
wire w2;    //: /sn:0 {0}(421,135)(615,135)(615,148)(625,148){1}
wire w5;    //: /sn:0 {0}(592,449)(738,449)(738,455)(766,455){1}
wire w9;    //: /sn:0 {0}(766,460)(613,460)(613,501)(603,501){1}
//: enddecls

  //: joint g44 (P12) @(184, 758) /w:[ 5 6 8 -1 ]
  or g4 (.I0(w2), .I1(G0), .Z(C4));   //: @(636,151) /sn:0 /delay:" 3" /w:[ 1 9 0 ]
  and g8 (.I0(C0), .I1(P0), .I2(P4), .Z(w3));   //: @(437,245) /sn:0 /delay:" 3" /w:[ 13 13 27 0 ]
  //: output g47 (C16) @(943,714) /sn:0 /w:[ 1 ]
  //: input g16 (G8) @(133,550) /sn:0 /w:[ 0 ]
  and g3 (.I0(P0), .I1(C0), .Z(w2));   //: @(411,135) /sn:0 /delay:" 3" /w:[ 9 0 0 ]
  //: joint g26 (G4) @(476, 331) /w:[ 6 -1 5 8 ]
  //: input g17 (P8) @(144,450) /sn:0 /w:[ 25 ]
  //: input g2 (P0) @(162,126) /sn:0 /w:[ 0 ]
  //: input g30 (G12) @(106,821) /sn:0 /w:[ 0 ]
  //: joint g23 (G0) @(237, 190) /w:[ 2 -1 1 16 ]
  //: joint g24 (P8) @(315, 450) /w:[ 6 -1 5 8 ]
  //: joint g39 (P12) @(143, 758) /w:[ 11 12 14 22 ]
  //: input g1 (G0) @(158,190) /sn:0 /w:[ 0 ]
  //: joint g60 (G4) @(391, 331) /w:[ 4 -1 3 10 ]
  //: output g29 (C12) @(919,465) /sn:0 /w:[ 0 ]
  //: joint g51 (P4) @(324, 289) /w:[ 2 -1 4 1 ]
  and g18 (.I0(C0), .I1(P0), .I2(P4), .I3(P8), .Z(w9));   //: @(593,501) /sn:0 /delay:" 3" /w:[ 11 17 19 7 1 ]
  and g25 (.I0(G4), .I1(P8), .Z(w6));   //: @(587,404) /sn:0 /delay:" 3" /w:[ 9 11 0 ]
  //: joint g10 (G0) @(291, 190) /w:[ 6 -1 5 12 ]
  or g65 (.I0(w0), .I1(G12), .I2(w16), .I3(w17), .Z(GG));   //: @(851,956) /sn:0 /delay:" 3" /w:[ 0 5 0 0 0 ]
  //: joint g64 (G0) @(322, 190) /w:[ 8 -1 7 10 ]
  and g49 (.I0(P0), .I1(P8), .I2(P4), .I3(P12), .Z(PG));   //: @(684,881) /sn:0 /delay:" 3" /w:[ 11 21 0 21 0 ]
  //: input g6 (P4) @(159,289) /sn:0 /w:[ 17 ]
  //: joint g50 (P0) @(365, 126) /w:[ 8 -1 7 10 ]
  //: joint g35 (P8) @(175, 450) /w:[ 13 14 16 28 ]
  //: joint g56 (G8) @(213, 553) /w:[ 2 -1 1 8 ]
  //: input g7 (G4) @(165,331) /sn:0 /w:[ 0 ]
  and g9 (.I0(G0), .I1(P4), .Z(w7));   //: @(422,281) /sn:0 /delay:" 3" /w:[ 13 3 0 ]
  //: joint g58 (P12) @(225, 758) /w:[ 2 -1 4 1 ]
  and g22 (.I0(G0), .I1(P4), .I2(P8), .Z(w5));   //: @(582,449) /sn:0 /delay:" 3" /w:[ 17 15 9 0 ]
  //: input g31 (P12) @(110,758) /sn:0 /w:[ 19 ]
  //: joint g59 (P8) @(208, 436) /w:[ 20 -1 19 22 ]
  //: output g67 (GG) @(963,957) /sn:0 /w:[ 1 ]
  //: joint g33 (P0) @(238, 126) /w:[ 4 -1 3 14 ]
  //: joint g45 (G8) @(431, 553) /w:[ 4 -1 3 6 ]
  and g54 (.I0(P12), .I1(G8), .Z(w0));   //: @(669,926) /sn:0 /delay:" 3" /w:[ 25 9 1 ]
  //: joint g41 (G4) @(292, 331) /w:[ 2 -1 1 12 ]
  and g36 (.I0(G0), .I1(P8), .I2(P4), .I3(P12), .Z(w10));   //: @(526,730) /sn:0 /delay:" 3" /w:[ 15 15 21 13 0 ]
  and g40 (.I0(G4), .I1(P8), .I2(P12), .Z(w11));   //: @(529,674) /sn:0 /delay:" 3" /w:[ 13 27 23 0 ]
  //: joint g42 (P8) @(159, 450) /w:[ 17 18 24 26 ]
  //: joint g52 (P12) @(125, 758) /w:[ 15 16 18 20 ]
  //: joint g66 (G12) @(260, 821) /w:[ 2 -1 1 4 ]
  //: joint g12 (C0) @(349, 137) /w:[ 1 -1 2 12 ]
  or g46 (.I0(w12), .I1(w11), .I2(w10), .I3(w4), .I4(G12), .Z(C16));   //: @(717,714) /sn:0 /delay:" 3" /w:[ 1 1 1 1 3 0 ]
  and g57 (.I0(G4), .I1(P8), .I2(P12), .Z(w16));   //: @(673,966) /sn:0 /delay:" 3" /w:[ 11 23 0 1 ]
  or g28 (.I0(w6), .I1(w5), .I2(w9), .I3(G8), .Z(C12));   //: @(777,457) /sn:0 /delay:" 3" /w:[ 1 1 0 5 1 ]
  //: joint g34 (P4) @(264, 289) /w:[ 9 -1 10 22 ]
  //: output g5 (C4) @(786,151) /sn:0 /w:[ 1 ]
  or g14 (.I0(w3), .I1(w7), .I2(G4), .Z(C8));   //: @(632,281) /sn:0 /delay:" 3" /w:[ 1 1 7 0 ]
  //: joint g11 (P0) @(307, 126) /w:[ 6 -1 5 12 ]
  //: joint g21 (P4) @(194, 289) /w:[ 13 14 16 18 ]
  //: joint g19 (C0) @(254, 137) /w:[ 3 -1 4 10 ]
  and g61 (.I0(G0), .I1(P4), .I2(P8), .I3(P12), .Z(w17));   //: @(681,1011) /sn:0 /delay:" 3" /w:[ 11 25 0 17 1 ]
  //: joint g20 (P0) @(216, 126) /w:[ 2 -1 1 16 ]
  and g32 (.I0(P0), .I1(C0), .I2(P4), .I3(P8), .I4(P12), .Z(w4));   //: @(526,773) /sn:0 /delay:" 3" /w:[ 15 9 23 29 3 0 ]
  //: joint g63 (P4) @(279, 289) /w:[ 7 -1 8 24 ]
  //: input g0 (C0) @(161,159) /sn:0 /w:[ 7 ]
  and g43 (.I0(G8), .I1(P12), .Z(w12));   //: @(521,603) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: output g15 (C8) @(796,282) /sn:0 /w:[ 1 ]
  //: joint g38 (P4) @(226, 289) /w:[ 11 -1 12 20 ]
  //: joint g48 (C0) @(198, 137) /w:[ 5 -1 6 8 ]
  //: joint g27 (P8) @(233, 450) /w:[ 4 10 3 -1 ]
  //: joint g62 (P8) @(201, 450) /w:[ 2 -1 12 1 ]
  //: joint g37 (G0) @(271, 190) /w:[ 4 -1 3 14 ]
  //: joint g55 (P12) @(168, 758) /w:[ 9 -1 10 24 ]
  //: output g53 (PG) @(953,881) /sn:0 /w:[ 1 ]
  //: joint g13 (P4) @(309, 289) /w:[ 5 -1 6 26 ]

endmodule

module CLA4BITS(C, COut, P, A, B, S, G);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] B;    //: /sn:0 {0}(124,-71)(124,23)(257,23){1}
//: {2}(258,23)(326,23){3}
//: {4}(327,23)(392,23){5}
//: {6}(393,23)(451,23){7}
//: {8}(452,23)(767,23){9}
input [3:0] A;    //: /sn:0 {0}(102,-69)(102,47)(238,47){1}
//: {2}(239,47)(307,47){3}
//: {4}(308,47)(367,47){5}
//: {6}(368,47)(429,47){7}
//: {8}(430,47)(790,47){9}
output G;    //: /sn:0 {0}(432,270)(432,355){1}
output P;    //: /sn:0 {0}(391,270)(391,314)(392,314)(392,341){1}
input C;    //: /sn:0 /dp:3 {0}(466,139)(521,139){1}
//: {2}(525,139)(557,139){3}
//: {4}(523,141)(523,254)(507,254){5}
output COut;    //: /sn:0 {0}(62,251)(176,251)(176,247)(190,247){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(46,186)(94,186){1}
wire w13;    //: /sn:0 {0}(341,135)(357,135)(357,228){1}
wire w16;    //: /sn:0 /dp:1 {0}(334,155)(334,191)(100,191){1}
wire w6;    //: /sn:0 {0}(258,27)(258,115){1}
wire w7;    //: /sn:0 {0}(239,51)(239,59)(241,59)(241,115){1}
wire w4;    //: /sn:0 {0}(308,51)(308,59)(309,59)(309,113){1}
wire w22;    //: /sn:0 {0}(404,138)(408,138)(408,162)(421,162)(421,207)(430,207)(430,228){1}
wire w3;    //: /sn:0 {0}(393,27)(393,114){1}
wire w0;    //: /sn:0 {0}(430,51)(430,59)(435,59)(435,116){1}
wire w20;    //: /sn:0 {0}(460,228)(460,214)(434,214)(434,158){1}
wire w12;    //: /sn:0 {0}(305,155)(305,218)(302,218)(302,228){1}
wire w18;    //: /sn:0 /dp:1 {0}(258,157)(258,201)(100,201){1}
wire w19;    //: /sn:0 {0}(248,157)(248,224)(253,224)(253,228){1}
wire w10;    //: /sn:0 {0}(458,158)(458,171)(100,171){1}
wire w23;    //: /sn:0 {0}(270,134)(287,134)(287,228){1}
wire w21;    //: /sn:0 {0}(487,228)(487,217)(463,217)(463,187)(445,187)(445,158){1}
wire w1;    //: /sn:0 {0}(452,27)(452,35)(455,35)(455,116){1}
wire w8;    //: /sn:0 {0}(367,228)(367,215)(370,215)(370,156){1}
wire w14;    //: /sn:0 {0}(394,156)(394,181)(100,181){1}
wire w2;    //: /sn:0 {0}(368,51)(368,59)(371,59)(371,114){1}
wire w11;    //: /sn:0 {0}(226,228)(226,180)(236,180)(236,157){1}
wire w15;    //: /sn:0 {0}(321,155)(321,228){1}
wire w5;    //: /sn:0 {0}(327,27)(327,35)(328,35)(328,113){1}
wire w9;    //: /sn:0 {0}(389,228)(389,200)(381,200)(381,156){1}
//: enddecls

  //: input g4 (C) @(559,139) /sn:0 /R:2 /w:[ 3 ]
  tran g8(.Z(w7), .I(A[3]));   //: @(239,45) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: joint g16 (C) @(523, 139) /w:[ 2 -1 1 4 ]
  PFA g3 (.B(w1), .A(w0), .C(C), .S(w10), .G(w21), .P(w20));   //: @(425, 117) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<1 ]
  //: output g17 (COut) @(65,251) /sn:0 /R:2 /w:[ 0 ]
  PFA g2 (.B(w3), .A(w2), .C(w22), .S(w14), .G(w9), .P(w8));   //: @(363, 115) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<1 Bo2<1 ]
  PFA g1 (.B(w5), .A(w4), .C(w13), .S(w16), .G(w15), .P(w12));   //: @(300, 114) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<0 Bo2<0 ]
  //: output g18 (P) @(392,338) /sn:0 /R:3 /w:[ 1 ]
  tran g10(.Z(w4), .I(A[2]));   //: @(308,45) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: input g6 (A) @(102,-71) /sn:0 /R:3 /w:[ 0 ]
  //: input g7 (B) @(124,-73) /sn:0 /R:3 /w:[ 0 ]
  tran g9(.Z(w6), .I(B[3]));   //: @(258,21) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g12(.Z(w2), .I(A[1]));   //: @(368,45) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  CLALogic g5 (.G3(w19), .P3(w11), .G2(w15), .P2(w12), .G1(w9), .P1(w8), .G0(w21), .P0(w20), .C0(C), .C3(w23), .C1(w22), .C2(w13), .C4(COut), .GG(G), .PG(P));   //: @(191, 229) /sz:(315, 40) /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Ti3>1 Ti4>0 Ti5>0 Ti6>0 Ti7>0 Ri0>5 To0<1 To1<1 To2<1 Lo0<1 Bo0<0 Bo1<0 ]
  tran g14(.Z(w0), .I(A[0]));   //: @(430,45) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g11(.Z(w5), .I(B[2]));   //: @(327,21) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: output g21 (S) @(49,186) /sn:0 /R:2 /w:[ 0 ]
  //: output g19 (G) @(432,352) /sn:0 /R:3 /w:[ 1 ]
  concat g20 (.I0(w10), .I1(w14), .I2(w16), .I3(w18), .Z(S));   //: @(95,186) /sn:0 /R:2 /w:[ 1 1 1 1 1 ] /dr:0
  PFA g0 (.B(w6), .A(w7), .C(w23), .S(w18), .G(w19), .P(w11));   //: @(229, 116) /sz:(40, 40) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>0 Bo0<0 Bo1<0 Bo2<1 ]
  tran g15(.Z(w1), .I(B[0]));   //: @(452,21) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g13(.Z(w3), .I(B[1]));   //: @(393,21) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1

endmodule

module CLALogic(C4, G2, P2, P0, G3, G0, C3, P1, G1, P3, GG, C1, C0, C2, PG);
//: interface  /sz:(40, 40) /bd:[ ]
input G2;    //: /sn:0 {0}(137,533)(191,533){1}
//: {2}(195,533)(409,533){3}
//: {4}(413,533)(738,533)(738,445)(746,445){5}
//: {6}(411,535)(411,580)(490,580){7}
//: {8}(193,535)(193,908)(638,908){9}
input C0;    //: /sn:0 /dp:3 {0}(380,117)(331,117){1}
//: {2}(327,117)(236,117){3}
//: {4}(232,117)(180,117){5}
//: {6}(176,117)(147,117)(147,139)(143,139){7}
//: {8}(178,119)(178,748)(495,748){9}
//: {10}(234,119)(234,474)(562,474){11}
//: {12}(329,119)(329,220)(406,220){13}
output GG;    //: /sn:0 /dp:1 {0}(841,935)(934,935)(934,937)(946,937){1}
input P1;    //: /sn:0 {0}(653,864)(304,864)(304,271){1}
//: {2}(306,269)(385,269)(385,263)(391,263){3}
//: {4}(302,269)(291,269){5}
//: {6}(287,269)(261,269){7}
//: {8}(257,269)(246,269){9}
//: {10}(242,269)(208,269){11}
//: {12}(204,269)(176,269){13}
//: {14}(174,267)(174,263)(152,263)(152,301)(197,301)(197,429)(551,429){15}
//: {16}(172,269)(141,269){17}
//: {18}(174,271)(174,484)(562,484){19}
//: {20}(206,271)(206,713)(495,713){21}
//: {22}(244,271)(244,753)(495,753){23}
//: {24}(259,271)(259,281)(267,281)(267,989)(649,989){25}
//: {26}(289,271)(289,339)(319,339)(319,230)(406,230){27}
output C3;    //: /sn:0 /dp:1 {0}(902,445)(848,445)(848,437)(767,437){1}
output PG;    //: /sn:0 {0}(674,861)(936,861){1}
input G0;    //: /sn:0 /dp:9 {0}(140,170)(215,170){1}
//: {2}(219,170)(249,170){3}
//: {4}(253,170)(269,170){5}
//: {6}(273,170)(300,170){7}
//: {8}(304,170)(647,170)(647,148)(599,148)(599,133)(605,133){9}
//: {10}(302,172)(302,984)(649,984){11}
//: {12}(271,172)(271,258)(391,258){13}
//: {14}(251,172)(251,703)(495,703){15}
//: {16}(217,172)(217,424)(551,424){17}
output C4;    //: /sn:0 {0}(707,694)(926,694){1}
output C2;    //: /sn:0 {0}(622,261)(769,261)(769,262)(779,262){1}
input P3;    //: /sn:0 {0}(642,951)(205,951)(205,740){1}
//: {2}(207,738)(259,738)(259,763)(495,763){3}
//: {4}(203,738)(166,738){5}
//: {6}(164,736)(164,585)(490,585){7}
//: {8}(162,738)(150,738){9}
//: {10}(146,738)(125,738){11}
//: {12}(123,736)(123,718)(495,718){13}
//: {14}(121,738)(107,738){15}
//: {16}(105,736)(105,726)(120,726)(120,999)(649,999){17}
//: {18}(103,738)(92,738){19}
//: {20}(105,740)(105,869)(653,869){21}
//: {22}(123,740)(123,750)(138,750)(138,659)(498,659){23}
//: {24}(148,740)(148,903)(638,903){25}
input G1;    //: /sn:0 /dp:11 {0}(147,311)(270,311){1}
//: {2}(274,311)(369,311){3}
//: {4}(373,311)(454,311){5}
//: {6}(458,311)(593,311)(593,266)(601,266){7}
//: {8}(456,313)(456,381)(556,381){9}
//: {10}(371,313)(371,941)(642,941){11}
//: {12}(272,313)(272,649)(498,649){13}
input G3;    //: /sn:0 {0}(88,801)(250,801){1}
//: {2}(254,801)(644,801)(644,704)(686,704){3}
//: {4}(252,803)(252,933)(820,933){5}
output C1;    //: /sn:0 {0}(626,131)(769,131){1}
input P0;    //: /sn:0 {0}(144,106)(194,106){1}
//: {2}(198,106)(216,106){3}
//: {4}(220,106)(285,106){5}
//: {6}(289,106)(343,106){7}
//: {8}(347,106)(374,106)(374,112)(380,112){9}
//: {10}(345,108)(345,854)(653,854){11}
//: {12}(287,108)(287,225)(406,225){13}
//: {14}(218,108)(218,743)(495,743){15}
//: {16}(196,108)(196,479)(562,479){17}
input P2;    //: /sn:0 /dp:21 {0}(649,994)(181,994)(181,432){1}
//: {2}(183,430)(211,430){3}
//: {4}(215,430)(293,430){5}
//: {6}(297,430)(355,430)(355,489)(562,489){7}
//: {8}(295,432)(295,466)(309,466)(309,434)(551,434){9}
//: {10}(213,428)(213,386)(556,386){11}
//: {12}(179,430)(157,430){13}
//: {14}(155,428)(155,418)(170,418)(170,708)(495,708){15}
//: {16}(153,430)(141,430){17}
//: {18}(139,428)(139,377)(159,377)(159,391)(170,391)(170,416)(186,416){19}
//: {20}(190,416)(292,416)(292,859)(653,859){21}
//: {22}(188,418)(188,946)(642,946){23}
//: {24}(137,430)(126,430){25}
//: {26}(139,432)(139,654)(498,654){27}
//: {28}(155,432)(155,758)(495,758){29}
wire w16;    //: /sn:0 {0}(820,938)(673,938)(673,946)(663,946){1}
wire w6;    //: /sn:0 {0}(577,384)(736,384)(736,430)(746,430){1}
wire w7;    //: /sn:0 {0}(412,261)(601,261){1}
wire w4;    //: /sn:0 {0}(516,753)(633,753)(633,699)(686,699){1}
wire w0;    //: /sn:0 /dp:1 {0}(820,928)(669,928)(669,906)(659,906){1}
wire w3;    //: /sn:0 {0}(427,225)(591,225)(591,256)(601,256){1}
wire w12;    //: /sn:0 {0}(511,583)(676,583)(676,684)(686,684){1}
wire w10;    //: /sn:0 {0}(516,710)(583,710)(583,694)(686,694){1}
wire w17;    //: /sn:0 {0}(820,943)(680,943)(680,991)(670,991){1}
wire w2;    //: /sn:0 {0}(401,115)(595,115)(595,128)(605,128){1}
wire w11;    //: /sn:0 {0}(519,654)(592,654)(592,681)(655,681)(655,689)(686,689){1}
wire w5;    //: /sn:0 {0}(572,429)(718,429)(718,435)(746,435){1}
wire w9;    //: /sn:0 {0}(746,440)(593,440)(593,481)(583,481){1}
//: enddecls

  //: joint g44 (P3) @(164, 738) /w:[ 5 6 8 -1 ]
  or g4 (.I0(w2), .I1(G0), .Z(C1));   //: @(616,131) /sn:0 /delay:" 3" /w:[ 1 9 0 ]
  and g8 (.I0(C0), .I1(P0), .I2(P1), .Z(w3));   //: @(417,225) /sn:0 /delay:" 3" /w:[ 13 13 27 0 ]
  //: output g47 (C4) @(923,694) /sn:0 /w:[ 1 ]
  //: input g16 (G2) @(135,533) /sn:0 /w:[ 0 ]
  and g3 (.I0(P0), .I1(C0), .Z(w2));   //: @(391,115) /sn:0 /delay:" 3" /w:[ 9 0 0 ]
  //: joint g26 (G1) @(456, 311) /w:[ 6 -1 5 8 ]
  //: input g17 (P2) @(124,430) /sn:0 /w:[ 25 ]
  //: input g2 (P0) @(142,106) /sn:0 /w:[ 0 ]
  //: input g30 (G3) @(86,801) /sn:0 /w:[ 0 ]
  //: joint g23 (G0) @(217, 170) /w:[ 2 -1 1 16 ]
  //: joint g24 (P2) @(295, 430) /w:[ 6 -1 5 8 ]
  //: joint g39 (P3) @(123, 738) /w:[ 11 12 14 22 ]
  //: input g1 (G0) @(138,170) /sn:0 /w:[ 0 ]
  //: joint g60 (G1) @(371, 311) /w:[ 4 -1 3 10 ]
  //: output g29 (C3) @(899,445) /sn:0 /w:[ 0 ]
  //: joint g51 (P1) @(304, 269) /w:[ 2 -1 4 1 ]
  and g18 (.I0(C0), .I1(P0), .I2(P1), .I3(P2), .Z(w9));   //: @(573,481) /sn:0 /delay:" 3" /w:[ 11 17 19 7 1 ]
  and g25 (.I0(G1), .I1(P2), .Z(w6));   //: @(567,384) /sn:0 /delay:" 3" /w:[ 9 11 0 ]
  //: joint g10 (G0) @(271, 170) /w:[ 6 -1 5 12 ]
  or g65 (.I0(w0), .I1(G3), .I2(w16), .I3(w17), .Z(GG));   //: @(831,935) /sn:0 /delay:" 3" /w:[ 0 5 0 0 0 ]
  //: joint g64 (G0) @(302, 170) /w:[ 8 -1 7 10 ]
  and g49 (.I0(P0), .I1(P2), .I2(P1), .I3(P3), .Z(PG));   //: @(664,861) /sn:0 /delay:" 3" /w:[ 11 21 0 21 0 ]
  //: input g6 (P1) @(139,269) /sn:0 /w:[ 17 ]
  //: joint g50 (P0) @(345, 106) /w:[ 8 -1 7 10 ]
  //: joint g35 (P2) @(155, 430) /w:[ 13 14 16 28 ]
  //: joint g56 (G2) @(193, 533) /w:[ 2 -1 1 8 ]
  //: input g7 (G1) @(145,311) /sn:0 /w:[ 0 ]
  and g9 (.I0(G0), .I1(P1), .Z(w7));   //: @(402,261) /sn:0 /delay:" 3" /w:[ 13 3 0 ]
  //: joint g58 (P3) @(205, 738) /w:[ 2 -1 4 1 ]
  and g22 (.I0(G0), .I1(P1), .I2(P2), .Z(w5));   //: @(562,429) /sn:0 /delay:" 3" /w:[ 17 15 9 0 ]
  //: input g31 (P3) @(90,738) /sn:0 /w:[ 19 ]
  //: joint g59 (P2) @(188, 416) /w:[ 20 -1 19 22 ]
  //: output g67 (GG) @(943,937) /sn:0 /w:[ 1 ]
  //: joint g33 (P0) @(218, 106) /w:[ 4 -1 3 14 ]
  //: joint g45 (G2) @(411, 533) /w:[ 4 -1 3 6 ]
  and g54 (.I0(P3), .I1(G2), .Z(w0));   //: @(649,906) /sn:0 /delay:" 3" /w:[ 25 9 1 ]
  //: joint g41 (G1) @(272, 311) /w:[ 2 -1 1 12 ]
  and g36 (.I0(G0), .I1(P2), .I2(P1), .I3(P3), .Z(w10));   //: @(506,710) /sn:0 /delay:" 3" /w:[ 15 15 21 13 0 ]
  and g40 (.I0(G1), .I1(P2), .I2(P3), .Z(w11));   //: @(509,654) /sn:0 /delay:" 3" /w:[ 13 27 23 0 ]
  //: joint g42 (P2) @(139, 430) /w:[ 17 18 24 26 ]
  //: joint g52 (P3) @(105, 738) /w:[ 15 16 18 20 ]
  //: joint g66 (G3) @(252, 801) /w:[ 2 -1 1 4 ]
  //: joint g12 (C0) @(329, 117) /w:[ 1 -1 2 12 ]
  or g46 (.I0(w12), .I1(w11), .I2(w10), .I3(w4), .I4(G3), .Z(C4));   //: @(697,694) /sn:0 /delay:" 3" /w:[ 1 1 1 1 3 0 ]
  and g57 (.I0(G1), .I1(P2), .I2(P3), .Z(w16));   //: @(653,946) /sn:0 /delay:" 3" /w:[ 11 23 0 1 ]
  or g28 (.I0(w6), .I1(w5), .I2(w9), .I3(G2), .Z(C3));   //: @(757,437) /sn:0 /delay:" 3" /w:[ 1 1 0 5 1 ]
  //: joint g34 (P1) @(244, 269) /w:[ 9 -1 10 22 ]
  //: output g5 (C1) @(766,131) /sn:0 /w:[ 1 ]
  or g14 (.I0(w3), .I1(w7), .I2(G1), .Z(C2));   //: @(612,261) /sn:0 /delay:" 3" /w:[ 1 1 7 0 ]
  //: joint g11 (P0) @(287, 106) /w:[ 6 -1 5 12 ]
  //: joint g21 (P1) @(174, 269) /w:[ 13 14 16 18 ]
  //: joint g19 (C0) @(234, 117) /w:[ 3 -1 4 10 ]
  and g61 (.I0(G0), .I1(P1), .I2(P2), .I3(P3), .Z(w17));   //: @(660,991) /sn:0 /delay:" 3" /w:[ 11 25 0 17 1 ]
  //: joint g20 (P0) @(196, 106) /w:[ 2 -1 1 16 ]
  and g32 (.I0(P0), .I1(C0), .I2(P1), .I3(P2), .I4(P3), .Z(w4));   //: @(506,753) /sn:0 /delay:" 3" /w:[ 15 9 23 29 3 0 ]
  //: joint g63 (P1) @(259, 269) /w:[ 7 -1 8 24 ]
  //: input g0 (C0) @(141,139) /sn:0 /w:[ 7 ]
  and g43 (.I0(G2), .I1(P3), .Z(w12));   //: @(501,583) /sn:0 /delay:" 3" /w:[ 7 7 0 ]
  //: output g15 (C2) @(776,262) /sn:0 /w:[ 1 ]
  //: joint g38 (P1) @(206, 269) /w:[ 11 -1 12 20 ]
  //: joint g48 (C0) @(178, 117) /w:[ 5 -1 6 8 ]
  //: joint g27 (P2) @(213, 430) /w:[ 4 10 3 -1 ]
  //: joint g62 (P2) @(181, 430) /w:[ 2 -1 12 1 ]
  //: joint g37 (G0) @(251, 170) /w:[ 4 -1 3 14 ]
  //: joint g55 (P3) @(148, 738) /w:[ 9 -1 10 24 ]
  //: output g53 (PG) @(933,861) /sn:0 /w:[ 1 ]
  //: joint g13 (P1) @(289, 269) /w:[ 5 -1 6 26 ]

endmodule

module main;    //: root_module
wire [15:0] w6;    //: /sn:0 {0}(525,199)(525,130)(535,130)(535,84){1}
wire w7;    //: /sn:0 {0}(239,325)(344,325)(344,322)(390,322){1}
wire w4;    //: /sn:0 {0}(232,234)(380,234)(380,227)(390,227){1}
wire [15:0] w0;    //: /sn:0 {0}(624,458)(624,507)(483,507)(483,365){1}
wire [15:0] w2;    //: /sn:0 /dp:1 {0}(438,199)(438,103)(394,103)(394,78){1}
wire w5;    //: /sn:0 {0}(239,277)(390,277){1}
wire w9;    //: /sn:0 {0}(579,291)(773,291){1}
//: enddecls

  //: dip g4 (w2) @(394,68) /sn:0 /w:[ 1 ] /st:10
  led g3 (.I(w5));   //: @(232,277) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: switch g2 (w9) @(791,291) /sn:0 /R:2 /w:[ 1 ] /st:1
  led g1 (.I(w0));   //: @(624,451) /sn:0 /w:[ 0 ] /type:3
  CLA16BITS g6 (.B(w6), .A(w2), .C(w9), .G(w4), .P(w7), .COut(w5), .S(w0));   //: @(391, 200) /sz:(187, 164) /sn:0 /p:[ Ti0>0 Ti1>0 Ri0>0 Lo0<1 Lo1<1 Lo2<1 Bo0<1 ]
  led g7 (.I(w7));   //: @(232,325) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: dip g5 (w6) @(535,74) /sn:0 /w:[ 1 ] /st:11
  led g0 (.I(w4));   //: @(225,234) /sn:0 /R:1 /w:[ 0 ] /type:0

endmodule
