//: version "1.8.7"

module CSA16(A, B, Cout, S, Cin);
//: interface  /sz:(40, 40) /bd:[ ]
input [15:0] B;    //: /sn:0 {0}(60,130)(238,130){1}
//: {2}(239,130)(484,130){3}
//: {4}(485,130)(712,130){5}
//: {6}(713,130)(949,130){7}
//: {8}(950,130)(1047,130){9}
input [15:0] A;    //: /sn:0 {0}(82,96)(183,96){1}
//: {2}(184,96)(412,96){3}
//: {4}(413,96)(654,96){5}
//: {6}(655,96)(892,96){7}
//: {8}(893,96)(1054,96){9}
output Cout;    //: /sn:0 {0}(64,257)(132,257)(132,263)(146,263){1}
input Cin;    //: /sn:0 {0}(1085,255)(1015,255){1}
output [15:0] S;    //: /sn:0 /dp:1 {0}(1020,433)(1074,433)(1074,432)(1084,432){1}
wire [3:0] w6;    //: /sn:0 {0}(655,100)(655,185){1}
wire [3:0] w7;    //: /sn:0 {0}(713,134)(713,137)(706,137)(706,185){1}
wire [3:0] w16;    //: /sn:0 {0}(239,134)(239,142)(235,142)(235,186){1}
wire w14;    //: /sn:0 {0}(381,266)(313,266)(313,268)(303,268){1}
wire [3:0] w19;    //: /sn:0 {0}(1014,418)(218,418)(218,340){1}
wire [3:0] w15;    //: /sn:0 {0}(184,100)(184,108)(183,108)(183,186){1}
wire w4;    //: /sn:0 {0}(849,266)(805,266)(805,264)(761,264){1}
wire [3:0] w3;    //: /sn:0 {0}(1014,448)(927,448)(927,340){1}
wire [3:0] w0;    //: /sn:0 {0}(893,100)(893,108)(894,108)(894,192){1}
wire [3:0] w1;    //: /sn:0 {0}(950,134)(950,142)(951,142)(951,192){1}
wire [3:0] w18;    //: /sn:0 {0}(1014,428)(455,428)(455,340){1}
wire [3:0] w12;    //: /sn:0 {0}(485,134)(485,143)(486,143)(486,191){1}
wire [3:0] w11;    //: /sn:0 {0}(413,100)(413,109)(421,109)(421,191){1}
wire [3:0] w5;    //: /sn:0 {0}(1014,438)(688,438)(688,338){1}
wire w9;    //: /sn:0 {0}(618,260)(552,260)(552,264)(541,264){1}
//: enddecls

  tran g8(.Z(w6), .I(A[7:4]));   //: @(655,94) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: input g4 (A) @(80,96) /sn:0 /w:[ 0 ]
  tran g13(.Z(w7), .I(B[7:4]));   //: @(713,128) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  CSA g3 (.B(w16), .A(w15), .C(w14), .COut(Cout), .S(w19));   //: @(147, 187) /sz:(155, 152) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<1 ]
  CSA g2 (.B(w12), .A(w11), .C(w9), .COut(w14), .S(w18));   //: @(382, 192) /sz:(158, 147) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  CPA g1 (.B(w1), .A(w0), .Cin(Cin), .Cout(w4), .S(w3));   //: @(850, 193) /sz:(164, 146) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  concat g16 (.I0(w3), .I1(w5), .I2(w18), .I3(w19), .Z(S));   //: @(1019,433) /sn:0 /w:[ 0 0 0 0 0 ] /dr:0
  tran g11(.Z(w16), .I(B[15:12]));   //: @(239,128) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g10(.Z(w1), .I(B[3:0]));   //: @(950,128) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g6(.Z(w15), .I(A[15:12]));   //: @(184,94) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g9 (B) @(58,130) /sn:0 /w:[ 0 ]
  tran g7(.Z(w11), .I(A[11:8]));   //: @(413,94) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: output g15 (Cout) @(67,257) /sn:0 /R:2 /w:[ 0 ]
  //: output g17 (S) @(1081,432) /sn:0 /w:[ 1 ]
  //: input g14 (Cin) @(1087,255) /sn:0 /R:2 /w:[ 0 ]
  tran g5(.Z(w0), .I(A[3:0]));   //: @(893,94) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  CSA g0 (.B(w7), .A(w6), .C(w4), .COut(w9), .S(w5));   //: @(619, 186) /sz:(141, 151) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  tran g12(.Z(w12), .I(B[11:8]));   //: @(485,128) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1

endmodule

module Full_Adder(COut, C, B, A, S);
//: interface  /sz:(40, 40) /bd:[ ]
input B;    //: /sn:0 /dp:1 {0}(240,107)(175,107){1}
//: {2}(171,107)(131,107)(131,151)(96,151){3}
//: {4}(173,109)(173,195)(317,195){5}
input A;    //: /sn:0 {0}(97,102)(142,102){1}
//: {2}(146,102)(240,102){3}
//: {4}(144,104)(144,200)(317,200){5}
output COut;    //: /sn:0 /dp:1 {0}(389,191)(422,191){1}
input C;    //: /sn:0 /dp:1 {0}(345,110)(295,110)(295,176){1}
//: {2}(297,178)(317,178){3}
//: {4}(295,180)(295,198)(95,198){5}
output S;    //: /sn:0 /dp:1 {0}(366,108)(389,108){1}
wire w0;    //: /sn:0 /dp:1 {0}(368,188)(344,188)(344,181)(338,181){1}
wire w1;    //: /sn:0 /dp:1 {0}(368,193)(345,193)(345,198)(338,198){1}
wire w2;    //: /sn:0 {0}(261,105)(274,105){1}
//: {2}(278,105)(345,105){3}
//: {4}(276,107)(276,183)(317,183){5}
//: enddecls

  and g8 (.I0(B), .I1(A), .Z(w1));   //: @(328,198) /sn:0 /delay:" 3" /w:[ 5 5 1 ]
  xor g4 (.I0(w2), .I1(C), .Z(S));   //: @(356,108) /sn:0 /delay:" 4" /w:[ 3 0 0 ]
  xor g3 (.I0(A), .I1(B), .Z(w2));   //: @(251,105) /sn:0 /delay:" 4" /w:[ 3 0 0 ]
  //: output g13 (COut) @(419,191) /sn:0 /w:[ 1 ]
  //: input g2 (C) @(93,198) /sn:0 /w:[ 5 ]
  //: input g1 (B) @(94,151) /sn:0 /w:[ 3 ]
  or g11 (.I0(w0), .I1(w1), .Z(COut));   //: @(379,191) /sn:0 /delay:" 3" /w:[ 0 0 0 ]
  //: joint g10 (A) @(144, 102) /w:[ 2 -1 1 4 ]
  //: joint g6 (w2) @(276, 105) /w:[ 2 -1 1 4 ]
  //: joint g9 (B) @(173, 107) /w:[ 1 -1 2 4 ]
  //: joint g7 (C) @(295, 178) /w:[ 2 1 -1 4 ]
  and g5 (.I0(C), .I1(w2), .Z(w0));   //: @(328,181) /sn:0 /delay:" 3" /w:[ 3 5 1 ]
  //: input g0 (A) @(95,102) /sn:0 /w:[ 0 ]
  //: output g12 (S) @(386,108) /sn:0 /w:[ 1 ]

endmodule

module CSA(B, C, S, A, COut);
//: interface  /sz:(40, 40) /bd:[ ]
supply1 w7;    //: /sn:0 /dp:1 {0}(355,160)(370,160){1}
input [3:0] B;    //: /sn:0 /dp:9 {0}(1,41)(85,41){1}
//: {2}(86,41)(159,41){3}
//: {4}(160,41)(222,41){5}
//: {6}(223,41)(282,41){7}
//: {8}(283,41)(323,41){9}
input [3:0] A;    //: /sn:0 /dp:9 {0}(53,25)(103,25){1}
//: {2}(104,25)(176,25){3}
//: {4}(177,25)(246,25){5}
//: {6}(247,25)(305,25){7}
//: {8}(306,25)(315,25){9}
output COut;    //: /sn:0 {0}(-35,157)(-46,157)(-46,118)(-56,118){1}
input C;    //: /sn:0 /dp:3 {0}(-45,318)(18,318){1}
//: {2}(22,318)(154,311)(154,312)(284,312){3}
//: {4}(20,316)(20,117)(-22,117)(-22,134){5}
supply1 w13;    //: /sn:0 {0}(372,98)(318,98){1}
output [3:0] S;    //: /sn:0 {0}(423,336)(307,336)(307,325){1}
wire w6;    //: /sn:0 {0}(215,185)(215,240)(113,240)(113,279){1}
wire S1;    //: /sn:0 {0}(83,180)(83,227)(133,227)(133,279){1}
wire C6;    //: /sn:0 {0}(109,170)(135,170){1}
wire w4;    //: /sn:0 {0}(156,182)(156,233)(123,233)(123,279){1}
wire C5;    //: /sn:0 {0}(177,169)(202,169){1}
wire A3;    //: /sn:0 {0}(104,29)(104,45){1}
//: {2}(102,47)(97,47)(97,66){3}
//: {4}(104,49)(104,138){5}
wire w0;    //: /sn:0 {0}(306,29)(306,52){1}
//: {2}(308,54)(314,54)(314,133){3}
//: {4}(306,56)(306,65){5}
wire w3;    //: /sn:0 {0}(103,279)(103,247)(285,247)(285,175){1}
wire A2;    //: /sn:0 {0}(177,29)(177,47)(169,47){1}
//: {2}(165,47)(161,47)(161,66){3}
//: {4}(167,49)(167,140){5}
wire B2;    //: /sn:0 {0}(160,45)(160,53)(156,53){1}
//: {2}(152,53)(146,53)(146,66){3}
//: {4}(154,55)(154,140){5}
wire C4;    //: /sn:0 {0}(276,168)(244,168){1}
wire C2;    //: /sn:0 {0}(177,96)(201,96){1}
wire w1;    //: /sn:0 {0}(283,45)(283,53){1}
//: {2}(285,55)(294,55)(294,133){3}
//: {4}(283,57)(283,65){5}
wire B1;    //: /sn:0 {0}(223,45)(223,55)(220,55){1}
//: {2}(216,55)(210,55)(210,66){3}
//: {4}(218,57)(218,143){5}
wire w18;    //: /sn:0 {0}(339,160)(318,160){1}
wire w8;    //: /sn:0 /dp:1 {0}(312,250)(312,219)(223,219)(223,108){1}
wire COut2;    //: /sn:0 {0}(135,99)(110,99){1}
wire COut1;    //: /sn:0 {0}(68,98)(4,98)(4,167)(-6,167){1}
wire w12;    //: /sn:0 {0}(-6,147)(28,147)(28,167)(64,167){1}
wire w2;    //: /sn:0 {0}(302,107)(302,250){1}
wire w11;    //: /sn:0 {0}(332,250)(332,213)(91,213)(91,109){1}
wire A1;    //: /sn:0 {0}(247,29)(247,47)(240,47){1}
//: {2}(236,47)(234,47)(234,66){3}
//: {4}(238,49)(238,143){5}
wire C1;    //: /sn:0 {0}(243,98)(274,98){1}
wire B3;    //: /sn:0 {0}(86,45)(86,53){1}
//: {2}(84,55)(77,55)(77,66){3}
//: {4}(86,57)(86,97)(75,97)(75,138){5}
wire [3:0] S3;    //: /sn:0 /dp:1 {0}(118,285)(118,286)(297,286)(297,296){1}
wire [3:0] w9;    //: /sn:0 /dp:1 {0}(317,256)(317,296){1}
wire S2;    //: /sn:0 /dp:1 {0}(162,108)(162,226)(322,226)(322,250){1}
//: enddecls

  tran g8(.Z(A2), .I(A[2]));   //: @(177,23) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  concat g4 (.I0(w2), .I1(w8), .I2(S2), .I3(w11), .Z(w9));   //: @(317,255) /sn:0 /R:3 /w:[ 1 0 1 0 0 ] /dr:0
  Full_Adder g3 (.B(B1), .A(A1), .C(C1), .COut(C2), .S(w8));   //: @(202, 67) /sz:(40, 40) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>0 Lo0<1 Bo0<1 ]
  concat g34 (.I0(w3), .I1(w6), .I2(w4), .I3(S1), .Z(S3));   //: @(118,284) /sn:0 /R:3 /w:[ 0 1 1 1 0 ] /dr:0
  not g37 (.I(w7), .Z(w18));   //: @(349,160) /sn:0 /R:2 /delay:" 4" /w:[ 0 0 ]
  tran g13(.Z(B1), .I(B[1]));   //: @(223,39) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  Full_Adder g2 (.B(w1), .A(w0), .C(w13), .COut(C1), .S(w2));   //: @(275, 66) /sz:(42, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Lo0<1 Bo0<0 ]
  Full_Adder g1 (.B(B2), .A(A2), .C(C2), .COut(COut2), .S(S2));   //: @(136, 67) /sz:(40, 40) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>0 Lo0<0 Bo0<0 ]
  mux g16 (.I0(S3), .I1(w9), .S(C), .Z(S));   //: @(307,312) /sn:0 /delay:" 2 2" /w:[ 1 1 3 1 ] /ss:0 /do:0
  tran g11(.Z(B3), .I(B[3]));   //: @(86,39) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: input g10 (B) @(-1,41) /sn:0 /w:[ 0 ]
  //: joint g28 (C) @(20, 318) /w:[ 2 4 1 -1 ]
  //: input g19 (C) @(-47,318) /sn:0 /w:[ 0 ]
  //: output g32 (S) @(420,336) /sn:0 /w:[ 0 ]
  //: joint g27 (B2) @(154, 53) /w:[ 1 -1 2 4 ]
  tran g6(.Z(w0), .I(A[0]));   //: @(306,23) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g9(.Z(A3), .I(A[3]));   //: @(104,23) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g7(.Z(A1), .I(A[1]));   //: @(247,23) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g31 (A3) @(104, 47) /w:[ -1 1 2 4 ]
  //: joint g20 (w1) @(283, 55) /w:[ 2 1 -1 4 ]
  //: supply1 g15 (w13) @(372,109) /sn:0 /R:3 /w:[ 0 ]
  mux g17 (.I0(w12), .I1(COut1), .S(C), .Z(COut));   //: @(-22,157) /sn:0 /R:3 /delay:" 2 2" /w:[ 0 1 5 0 ] /ss:0 /do:0
  Full_Adder g29 (.B(B3), .A(A3), .C(C6), .COut(w12), .S(S1));   //: @(65, 139) /sz:(43, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<1 Bo0<0 ]
  Full_Adder g25 (.B(B2), .A(A2), .C(C5), .COut(C6), .S(w4));   //: @(136, 141) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>0 Lo0<1 Bo0<0 ]
  tran g14(.Z(w1), .I(B[0]));   //: @(283,39) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  //: input g5 (A) @(51,25) /sn:0 /w:[ 0 ]
  //: joint g24 (A1) @(238, 47) /w:[ 1 -1 2 4 ]
  //: supply1 g36 (w7) @(370,171) /sn:0 /R:3 /w:[ 1 ]
  //: joint g21 (w0) @(306, 54) /w:[ 2 1 -1 4 ]
  //: joint g23 (B1) @(218, 55) /w:[ 1 -1 2 4 ]
  //: joint g26 (A2) @(167, 47) /w:[ 1 -1 2 4 ]
  Full_Adder g22 (.A(A1), .B(B1), .C(C4), .COut(C5), .S(w6));   //: @(203, 144) /sz:(40, 40) /sn:0 /p:[ Ti0>5 Ti1>5 Ri0>1 Lo0<1 Bo0<0 ]
  Full_Adder g0 (.A(A3), .B(B3), .C(COut2), .COut(COut1), .S(w11));   //: @(69, 67) /sz:(40, 41) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>1 Lo0<0 Bo0<1 ]
  Full_Adder g18 (.B(w1), .A(w0), .C(w18), .COut(C4), .S(w3));   //: @(277, 134) /sz:(40, 40) /sn:0 /p:[ Ti0>3 Ti1>3 Ri0>1 Lo0<0 Bo0<1 ]
  tran g12(.Z(B2), .I(B[2]));   //: @(160,39) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: joint g30 (B3) @(86, 55) /w:[ -1 1 2 4 ]
  //: output g33 (COut) @(-53,118) /sn:0 /R:2 /w:[ 1 ]

endmodule

module CPA(Cin, B, A, S, Cout);
//: interface  /sz:(40, 40) /bd:[ ]
input [3:0] B;    //: /sn:0 {0}(120,139)(325,139){1}
//: {2}(326,139)(552,139){3}
//: {4}(553,139)(743,139){5}
//: {6}(744,139)(945,139){7}
//: {8}(946,139)(1053,139){9}
input [3:0] A;    //: /sn:0 {0}(148,106)(287,106){1}
//: {2}(288,106)(499,106){3}
//: {4}(500,106)(709,106){5}
//: {6}(710,106)(905,106){7}
//: {8}(906,106)(1053,106){9}
output Cout;    //: /sn:0 {0}(153,249)(199,249)(199,248)(244,248){1}
input Cin;    //: /sn:0 {0}(1089,243)(1000,243){1}
output [3:0] S;    //: /sn:0 /dp:1 {0}(603,427)(603,465)(653,465){1}
wire w6;    //: /sn:0 {0}(553,143)(553,151)(551,151)(551,180){1}
wire w16;    //: /sn:0 {0}(946,143)(946,151)(949,151)(949,175){1}
wire w14;    //: /sn:0 {0}(669,251)(607,251)(607,245)(597,245){1}
wire w19;    //: /sn:0 {0}(877,243)(810,243){1}
wire w15;    //: /sn:0 {0}(906,110)(906,118)(905,118)(905,175){1}
wire w3;    //: /sn:0 /dp:1 {0}(298,309)(298,348)(618,348)(618,421){1}
wire w0;    //: /sn:0 {0}(288,110)(288,118)(286,118)(286,180){1}
wire w1;    //: /sn:0 {0}(326,143)(326,151)(327,151)(327,180){1}
wire w18;    //: /sn:0 {0}(931,311)(931,339)(588,339)(588,421){1}
wire w12;    //: /sn:0 {0}(608,421)(608,324)(542,324)(542,313){1}
wire w11;    //: /sn:0 {0}(744,143)(744,151)(747,151)(747,179){1}
wire w10;    //: /sn:0 {0}(710,110)(710,118)(709,118)(709,179){1}
wire w13;    //: /sn:0 {0}(738,311)(738,364)(598,364)(598,421){1}
wire w5;    //: /sn:0 {0}(500,110)(500,180){1}
wire w9;    //: /sn:0 {0}(462,252)(384,252)(384,235)(374,235){1}
//: enddecls

  tran g8(.Z(w10), .I(A[1]));   //: @(710,104) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: input g4 (Cin) @(1091,243) /sn:0 /R:2 /w:[ 0 ]
  tran g13(.Z(w1), .I(B[3]));   //: @(326,137) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  Full_Adder g3 (.B(w16), .A(w15), .C(Cin), .COut(w19), .S(w18));   //: @(878, 176) /sz:(121, 134) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  Full_Adder g2 (.B(w11), .A(w10), .C(w19), .COut(w14), .S(w13));   //: @(670, 180) /sz:(139, 130) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<0 ]
  Full_Adder g1 (.B(w6), .A(w5), .C(w14), .COut(w9), .S(w12));   //: @(463, 181) /sz:(133, 131) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<0 Bo0<1 ]
  concat g16 (.I0(w18), .I1(w13), .I2(w12), .I3(w3), .Z(S));   //: @(603,426) /sn:0 /R:3 /w:[ 1 1 0 1 0 ] /dr:0
  //: input g11 (B) @(118,139) /sn:0 /w:[ 0 ]
  tran g10(.Z(w5), .I(A[2]));   //: @(500,104) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: input g6 (A) @(146,106) /sn:0 /w:[ 0 ]
  tran g9(.Z(w0), .I(A[3]));   //: @(288,104) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  tran g7(.Z(w15), .I(A[0]));   //: @(906,104) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  tran g15(.Z(w11), .I(B[1]));   //: @(744,137) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: output g17 (S) @(650,465) /sn:0 /w:[ 1 ]
  tran g14(.Z(w6), .I(B[2]));   //: @(553,137) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  //: output g5 (Cout) @(156,249) /sn:0 /R:2 /w:[ 0 ]
  Full_Adder g0 (.B(w1), .A(w0), .C(w9), .COut(Cout), .S(w3));   //: @(245, 181) /sz:(128, 127) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]
  tran g12(.Z(w16), .I(B[0]));   //: @(946,137) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1

endmodule

module main;    //: root_module
wire [15:0] w4;    //: /sn:0 {0}(84,-82)(84,-32)(83,-32)(83,-23){1}
wire [15:0] w0;    //: /sn:0 {0}(163,270)(163,346)(263,346)(263,321){1}
wire [15:0] w1;    //: /sn:0 {0}(223,-80)(223,-23){1}
wire w2;    //: /sn:0 {0}(383,87)(383,119)(339,119){1}
wire w5;    //: /sn:0 {0}(-57,81)(-57,115)(-6,115){1}
//: enddecls

  //: switch g4 (w2) @(383,74) /sn:0 /R:3 /w:[ 0 ] /st:0
  //: dip g3 (w1) @(223,-90) /sn:0 /w:[ 0 ] /st:0
  //: dip g2 (w4) @(84,-92) /sn:0 /w:[ 0 ] /st:0
  led g1 (.I(w5));   //: @(-57,74) /sn:0 /w:[ 0 ] /type:0
  led g5 (.I(w0));   //: @(263,314) /sn:0 /w:[ 1 ] /type:3
  CSA16 g0 (.B(w1), .A(w4), .Cin(w2), .Cout(w5), .S(w0));   //: @(-5, -22) /sz:(343, 291) /sn:0 /p:[ Ti0>1 Ti1>1 Ri0>1 Lo0<1 Bo0<0 ]

endmodule
