//: version "1.8.7"

module HA(s, b, a, c);
//: interface  /sz:(166, 122) /bd:[ Ti0>b(113/166) Ti1>a(50/166) Lo0<c(59/122) Bo0<s(80/166) ]
input b;    //: /sn:0 {0}(259,188)(281,188){1}
//: {2}(285,188)(321,188)(321,179)(329,179){3}
//: {4}(283,190)(283,235)(330,235){5}
output s;    //: /sn:0 /dp:1 {0}(350,177)(426,177){1}
input a;    //: /sn:0 {0}(260,174)(295,174){1}
//: {2}(299,174)(329,174){3}
//: {4}(297,176)(297,230)(330,230){5}
output c;    //: /sn:0 /dp:1 {0}(351,233)(423,233){1}
//: enddecls

  //: output g4 (s) @(423,177) /sn:0 /w:[ 1 ]
  //: input g3 (b) @(257,188) /sn:0 /w:[ 0 ]
  //: input g2 (a) @(258,174) /sn:0 /w:[ 0 ]
  and g1 (.I0(a), .I1(b), .Z(c));   //: @(341,233) /sn:0 /delay:" 3" /w:[ 5 5 0 ]
  //: joint g6 (a) @(297, 174) /w:[ 2 -1 1 4 ]
  //: joint g7 (b) @(283, 188) /w:[ 2 -1 1 4 ]
  //: output g5 (c) @(420,233) /sn:0 /w:[ 1 ]
  xor g0 (.I0(a), .I1(b), .Z(s));   //: @(340,177) /sn:0 /delay:" 4" /w:[ 3 3 0 ]

endmodule

module main;    //: root_module
wire w4;    //: /sn:0 {0}(407,112)(414,112)(414,163){1}
wire w3;    //: /sn:0 /dp:1 {0}(265,255)(265,275)(332,275){1}
wire w0;    //: /sn:0 /dp:1 {0}(437,443)(437,453)(462,453)(462,396){1}
wire w1;    //: /sn:0 {0}(500,115)(516,115)(516,163){1}
//: enddecls

  led g4 (.I(w3));   //: @(265,248) /sn:0 /w:[ 0 ] /type:0
  led g3 (.I(w0));   //: @(437,436) /sn:0 /w:[ 0 ] /type:0
  //: switch g2 (w1) @(483,115) /sn:0 /w:[ 0 ] /st:0
  //: switch g1 (w4) @(390,112) /sn:0 /w:[ 0 ] /st:0
  HA g0 (.a(w4), .b(w1), .c(w3), .s(w0));   //: @(333, 164) /sz:(269, 231) /sn:0 /p:[ Ti0>1 Ti1>1 Lo0<1 Bo0<1 ]

endmodule
